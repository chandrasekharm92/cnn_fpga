`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:08:09 11/08/2017 
// Design Name: 
// Module Name:    cnn 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module cnn(weight1l0,weight1l1,weight1l2,weight1l3,weight1l4,weight1l5,weight1l6,weight1l7,weight1l8,weight1l9,weight1l10,weight1l11,weight1l12,weight1l13,weight1l14,weight1l15,weight1l16,weight1l17,weight1l18,weight1l19,weight1l20,weight1l21,weight1l22,weight1l23,weight1l24,
weight2l0,weight2l1,weight2l2,weight2l3,weight2l4,weight2l5,weight2l6,weight2l7,weight2l8,weight2l9,weight2l10,weight2l11,weight2l12,weight2l13,weight2l14,weight2l15,weight2l16,weight2l17,weight2l18,weight2l19,weight2l20,weight2l21,weight2l22,weight2l23,weight2l24,weight2l25,weight2l26,weight2l27,weight2l28,weight2l29,weight2l30,weight2l31,weight2l32,weight2l33,weight2l34,weight2l35,weight2l36,weight2l37,weight2l38,weight2l39,weight2l40,weight2l41,weight2l42,weight2l43,weight2l44,weight2l45,weight2l46,weight2l47,weight2l48,weight2l49,weight2l50,weight2l51,weight2l52,weight2l53,weight2l54,weight2l55,weight2l56,weight2l57,weight2l58,weight2l59,weight2l60,weight2l61,weight2l62,weight2l63,weight2l64,weight2l65,weight2l66,weight2l67,weight2l68,weight2l69,weight2l70,weight2l71,weight2l72,weight2l73,weight2l74,weight2l75,weight2l76,weight2l77,weight2l78,weight2l79,weight2l80,weight2l81,weight2l82,weight2l83,weight2l84,weight2l85,weight2l86,weight2l87,weight2l88,weight2l89,weight2l90,weight2l91,weight2l92,weight2l93,weight2l94,weight2l95,weight2l96,weight2l97,weight2l98,weight2l99,weight2l100,weight2l101,weight2l102,weight2l103,weight2l104,weight2l105,weight2l106,weight2l107,weight2l108,weight2l109,weight2l110,weight2l111,weight2l112,weight2l113,weight2l114,weight2l115,weight2l116,weight2l117,weight2l118,weight2l119,weight2l120,weight2l121,weight2l122,weight2l123,weight2l124,weight2l125,weight2l126,weight2l127,weight2l128,weight2l129,weight2l130,weight2l131,weight2l132,weight2l133,weight2l134,weight2l135,weight2l136,weight2l137,weight2l138,weight2l139,weight2l140,weight2l141,weight2l142,weight2l143,
in0,in1,in2,in3,in4,in5,in6,in7,in8,in9,in10,in11,in12,in13,in14,in15,in16,in17,in18,in19,in20,in21,in22,in23,in24,in25,in26,in27,in28,in29,in30,in31,in32,in33,in34,in35,in36,in37,in38,in39,in40,in41,in42,in43,in44,in45,in46,in47,in48,in49,in50,in51,in52,in53,in54,in55,in56,in57,in58,in59,in60,in61,in62,in63,in64,in65,in66,in67,in68,in69,in70,in71,in72,in73,in74,in75,in76,in77,in78,in79,in80,in81,in82,in83,in84,in85,in86,in87,in88,in89,in90,in91,in92,in93,in94,in95,in96,in97,in98,in99,in100,in101,in102,in103,in104,in105,in106,in107,in108,in109,in110,in111,in112,in113,in114,in115,in116,in117,in118,in119,in120,in121,in122,in123,in124,in125,in126,in127,in128,in129,in130,in131,in132,in133,in134,in135,in136,in137,in138,in139,in140,in141,in142,in143,in144,in145,in146,in147,in148,in149,in150,in151,in152,in153,in154,in155,in156,in157,in158,in159,in160,in161,in162,in163,in164,in165,in166,in167,in168,in169,in170,in171,in172,in173,in174,in175,in176,in177,in178,in179,in180,in181,in182,in183,in184,in185,in186,in187,in188,in189,in190,in191,in192,in193,in194,in195,in196,in197,in198,in199,in200,in201,in202,in203,in204,in205,in206,in207,in208,in209,in210,in211,in212,in213,in214,in215,in216,in217,in218,in219,in220,in221,in222,in223,in224,in225,in226,in227,in228,in229,in230,in231,in232,in233,in234,in235,in236,in237,in238,in239,in240,in241,in242,in243,in244,in245,in246,in247,in248,in249,in250,in251,in252,in253,in254,in255,in256,in257,in258,in259,in260,in261,in262,in263,in264,in265,in266,in267,in268,in269,in270,in271,in272,in273,in274,in275,in276,in277,in278,in279,in280,in281,in282,in283,in284,in285,in286,in287,in288,in289,in290,in291,in292,in293,in294,in295,in296,in297,in298,in299,in300,in301,in302,in303,in304,in305,in306,in307,in308,in309,in310,in311,in312,in313,in314,in315,in316,in317,in318,in319,in320,in321,in322,in323,in324,in325,in326,in327,in328,in329,in330,in331,in332,in333,in334,in335,in336,in337,in338,in339,in340,in341,in342,in343,in344,in345,in346,in347,in348,in349,in350,in351,in352,in353,in354,in355,in356,in357,in358,in359,in360,in361,in362,in363,in364,in365,in366,in367,in368,in369,in370,in371,in372,in373,in374,in375,in376,in377,in378,in379,in380,in381,in382,in383,in384,in385,in386,in387,in388,in389,in390,in391,in392,in393,in394,in395,in396,in397,in398,in399,in400,in401,in402,in403,in404,in405,in406,in407,in408,in409,in410,in411,in412,in413,in414,in415,in416,in417,in418,in419,in420,in421,in422,in423,in424,in425,in426,in427,in428,in429,in430,in431,in432,in433,in434,in435,in436,in437,in438,in439,in440,in441,in442,in443,in444,in445,in446,in447,in448,in449,in450,in451,in452,in453,in454,in455,in456,in457,in458,in459,in460,in461,in462,in463,in464,in465,in466,in467,in468,in469,in470,in471,in472,in473,in474,in475,in476,in477,in478,in479,in480,in481,in482,in483,in484,in485,in486,in487,in488,in489,in490,in491,in492,in493,in494,in495,in496,in497,in498,in499,in500,in501,in502,in503,in504,in505,in506,in507,in508,in509,in510,in511,in512,in513,in514,in515,in516,in517,in518,in519,in520,in521,in522,in523,in524,in525,in526,in527,in528,in529,in530,in531,in532,in533,in534,in535,in536,in537,in538,in539,in540,in541,in542,in543,in544,in545,in546,in547,in548,in549,in550,in551,in552,in553,in554,in555,in556,in557,in558,in559,in560,in561,in562,in563,in564,in565,in566,in567,in568,in569,in570,in571,in572,in573,in574,in575,in576,in577,in578,in579,in580,in581,in582,in583,in584,in585,in586,in587,in588,in589,in590,in591,in592,in593,in594,in595,in596,in597,in598,in599,in600,in601,in602,in603,in604,in605,in606,in607,in608,in609,in610,in611,in612,in613,in614,in615,in616,in617,in618,in619,in620,in621,in622,in623,in624,in625,in626,in627,in628,in629,in630,in631,in632,in633,in634,in635,in636,in637,in638,in639,in640,in641,in642,in643,in644,in645,in646,in647,in648,in649,in650,in651,in652,in653,in654,in655,in656,in657,in658,in659,in660,in661,in662,in663,in664,in665,in666,in667,in668,in669,in670,in671,in672,in673,in674,in675,in676,in677,in678,in679,in680,in681,in682,in683,in684,in685,in686,in687,in688,in689,in690,in691,in692,in693,in694,in695,in696,in697,in698,in699,in700,in701,in702,in703,in704,in705,in706,in707,in708,in709,in710,in711,in712,in713,in714,in715,in716,in717,in718,in719,in720,in721,in722,in723,in724,in725,in726,in727,in728,in729,in730,in731,in732,in733,in734,in735,in736,in737,in738,in739,in740,in741,in742,in743,in744,in745,in746,in747,in748,in749,in750,in751,in752,in753,in754,in755,in756,in757,in758,in759,in760,in761,in762,in763,in764,in765,in766,in767,in768,in769,in770,in771,in772,in773,in774,in775,in776,in777,in778,in779,in780,in781,in782,in783,
bias,clk,start,ready,out);

input [7:0] weight1l0;input [7:0] weight1l1;input [7:0] weight1l2;input [7:0] weight1l3;input [7:0] weight1l4;input [7:0] weight1l5;input [7:0] weight1l6;input [7:0] weight1l7;input [7:0] weight1l8;input [7:0] weight1l9;input [7:0] weight1l10;input [7:0] weight1l11;input [7:0] weight1l12;input [7:0] weight1l13;input [7:0] weight1l14;input [7:0] weight1l15;input [7:0] weight1l16;input [7:0] weight1l17;input [7:0] weight1l18;input [7:0] weight1l19;input [7:0] weight1l20;input [7:0] weight1l21;input [7:0] weight1l22;input [7:0] weight1l23;input [7:0] weight1l24;
input [7:0] weight2l0;input [7:0] weight2l1;input [7:0] weight2l2;input [7:0] weight2l3;input [7:0] weight2l4;input [7:0] weight2l5;input [7:0] weight2l6;input [7:0] weight2l7;input [7:0] weight2l8;input [7:0] weight2l9;input [7:0] weight2l10;input [7:0] weight2l11;input [7:0] weight2l12;input [7:0] weight2l13;input [7:0] weight2l14;input [7:0] weight2l15;input [7:0] weight2l16;input [7:0] weight2l17;input [7:0] weight2l18;input [7:0] weight2l19;input [7:0] weight2l20;input [7:0] weight2l21;input [7:0] weight2l22;input [7:0] weight2l23;input [7:0] weight2l24;input [7:0] weight2l25;input [7:0] weight2l26;input [7:0] weight2l27;input [7:0] weight2l28;input [7:0] weight2l29;input [7:0] weight2l30;input [7:0] weight2l31;input [7:0] weight2l32;input [7:0] weight2l33;input [7:0] weight2l34;input [7:0] weight2l35;input [7:0] weight2l36;input [7:0] weight2l37;input [7:0] weight2l38;input [7:0] weight2l39;input [7:0] weight2l40;input [7:0] weight2l41;input [7:0] weight2l42;input [7:0] weight2l43;input [7:0] weight2l44;input [7:0] weight2l45;input [7:0] weight2l46;input [7:0] weight2l47;input [7:0] weight2l48;input [7:0] weight2l49;input [7:0] weight2l50;input [7:0] weight2l51;input [7:0] weight2l52;input [7:0] weight2l53;input [7:0] weight2l54;input [7:0] weight2l55;input [7:0] weight2l56;input [7:0] weight2l57;input [7:0] weight2l58;input [7:0] weight2l59;input [7:0] weight2l60;input [7:0] weight2l61;input [7:0] weight2l62;input [7:0] weight2l63;input [7:0] weight2l64;input [7:0] weight2l65;input [7:0] weight2l66;input [7:0] weight2l67;input [7:0] weight2l68;input [7:0] weight2l69;input [7:0] weight2l70;input [7:0] weight2l71;input [7:0] weight2l72;input [7:0] weight2l73;input [7:0] weight2l74;input [7:0] weight2l75;input [7:0] weight2l76;input [7:0] weight2l77;input [7:0] weight2l78;input [7:0] weight2l79;input [7:0] weight2l80;input [7:0] weight2l81;input [7:0] weight2l82;input [7:0] weight2l83;input [7:0] weight2l84;input [7:0] weight2l85;input [7:0] weight2l86;input [7:0] weight2l87;input [7:0] weight2l88;input [7:0] weight2l89;input [7:0] weight2l90;input [7:0] weight2l91;input [7:0] weight2l92;input [7:0] weight2l93;input [7:0] weight2l94;input [7:0] weight2l95;input [7:0] weight2l96;input [7:0] weight2l97;input [7:0] weight2l98;input [7:0] weight2l99;input [7:0] weight2l100;input [7:0] weight2l101;input [7:0] weight2l102;input [7:0] weight2l103;input [7:0] weight2l104;input [7:0] weight2l105;input [7:0] weight2l106;input [7:0] weight2l107;input [7:0] weight2l108;input [7:0] weight2l109;input [7:0] weight2l110;input [7:0] weight2l111;input [7:0] weight2l112;input [7:0] weight2l113;input [7:0] weight2l114;input [7:0] weight2l115;input [7:0] weight2l116;input [7:0] weight2l117;input [7:0] weight2l118;input [7:0] weight2l119;input [7:0] weight2l120;input [7:0] weight2l121;input [7:0] weight2l122;input [7:0] weight2l123;input [7:0] weight2l124;input [7:0] weight2l125;input [7:0] weight2l126;input [7:0] weight2l127;input [7:0] weight2l128;input [7:0] weight2l129;input [7:0] weight2l130;input [7:0] weight2l131;input [7:0] weight2l132;input [7:0] weight2l133;input [7:0] weight2l134;input [7:0] weight2l135;input [7:0] weight2l136;input [7:0] weight2l137;input [7:0] weight2l138;input [7:0] weight2l139;input [7:0] weight2l140;input [7:0] weight2l141;input [7:0] weight2l142;input [7:0] weight2l143;
input [7:0] in0;input [7:0] in1;input [7:0] in2;input [7:0] in3;input [7:0] in4;input [7:0] in5;input [7:0] in6;input [7:0] in7;input [7:0] in8;input [7:0] in9;input [7:0] in10;input [7:0] in11;input [7:0] in12;input [7:0] in13;input [7:0] in14;input [7:0] in15;input [7:0] in16;input [7:0] in17;input [7:0] in18;input [7:0] in19;input [7:0] in20;input [7:0] in21;input [7:0] in22;input [7:0] in23;input [7:0] in24;input [7:0] in25;input [7:0] in26;input [7:0] in27;input [7:0] in28;input [7:0] in29;input [7:0] in30;input [7:0] in31;input [7:0] in32;input [7:0] in33;input [7:0] in34;input [7:0] in35;input [7:0] in36;input [7:0] in37;input [7:0] in38;input [7:0] in39;input [7:0] in40;input [7:0] in41;input [7:0] in42;input [7:0] in43;input [7:0] in44;input [7:0] in45;input [7:0] in46;input [7:0] in47;input [7:0] in48;input [7:0] in49;input [7:0] in50;input [7:0] in51;input [7:0] in52;input [7:0] in53;input [7:0] in54;input [7:0] in55;input [7:0] in56;input [7:0] in57;input [7:0] in58;input [7:0] in59;input [7:0] in60;input [7:0] in61;input [7:0] in62;input [7:0] in63;input [7:0] in64;input [7:0] in65;input [7:0] in66;input [7:0] in67;input [7:0] in68;input [7:0] in69;input [7:0] in70;input [7:0] in71;input [7:0] in72;input [7:0] in73;input [7:0] in74;input [7:0] in75;input [7:0] in76;input [7:0] in77;input [7:0] in78;input [7:0] in79;input [7:0] in80;input [7:0] in81;input [7:0] in82;input [7:0] in83;input [7:0] in84;input [7:0] in85;input [7:0] in86;input [7:0] in87;input [7:0] in88;input [7:0] in89;input [7:0] in90;input [7:0] in91;input [7:0] in92;input [7:0] in93;input [7:0] in94;input [7:0] in95;input [7:0] in96;input [7:0] in97;input [7:0] in98;input [7:0] in99;input [7:0] in100;input [7:0] in101;input [7:0] in102;input [7:0] in103;input [7:0] in104;input [7:0] in105;input [7:0] in106;input [7:0] in107;input [7:0] in108;input [7:0] in109;input [7:0] in110;input [7:0] in111;input [7:0] in112;input [7:0] in113;input [7:0] in114;input [7:0] in115;input [7:0] in116;input [7:0] in117;input [7:0] in118;input [7:0] in119;input [7:0] in120;input [7:0] in121;input [7:0] in122;input [7:0] in123;input [7:0] in124;input [7:0] in125;input [7:0] in126;input [7:0] in127;input [7:0] in128;input [7:0] in129;input [7:0] in130;input [7:0] in131;input [7:0] in132;input [7:0] in133;input [7:0] in134;input [7:0] in135;input [7:0] in136;input [7:0] in137;input [7:0] in138;input [7:0] in139;input [7:0] in140;input [7:0] in141;input [7:0] in142;input [7:0] in143;input [7:0] in144;input [7:0] in145;input [7:0] in146;input [7:0] in147;input [7:0] in148;input [7:0] in149;input [7:0] in150;input [7:0] in151;input [7:0] in152;input [7:0] in153;input [7:0] in154;input [7:0] in155;input [7:0] in156;input [7:0] in157;input [7:0] in158;input [7:0] in159;input [7:0] in160;input [7:0] in161;input [7:0] in162;input [7:0] in163;input [7:0] in164;input [7:0] in165;input [7:0] in166;input [7:0] in167;input [7:0] in168;input [7:0] in169;input [7:0] in170;input [7:0] in171;input [7:0] in172;input [7:0] in173;input [7:0] in174;input [7:0] in175;input [7:0] in176;input [7:0] in177;input [7:0] in178;input [7:0] in179;input [7:0] in180;input [7:0] in181;input [7:0] in182;input [7:0] in183;input [7:0] in184;input [7:0] in185;input [7:0] in186;input [7:0] in187;input [7:0] in188;input [7:0] in189;input [7:0] in190;input [7:0] in191;input [7:0] in192;input [7:0] in193;input [7:0] in194;input [7:0] in195;input [7:0] in196;input [7:0] in197;input [7:0] in198;input [7:0] in199;input [7:0] in200;input [7:0] in201;input [7:0] in202;input [7:0] in203;input [7:0] in204;input [7:0] in205;input [7:0] in206;input [7:0] in207;input [7:0] in208;input [7:0] in209;input [7:0] in210;input [7:0] in211;input [7:0] in212;input [7:0] in213;input [7:0] in214;input [7:0] in215;input [7:0] in216;input [7:0] in217;input [7:0] in218;input [7:0] in219;input [7:0] in220;input [7:0] in221;input [7:0] in222;input [7:0] in223;input [7:0] in224;input [7:0] in225;input [7:0] in226;input [7:0] in227;input [7:0] in228;input [7:0] in229;input [7:0] in230;input [7:0] in231;input [7:0] in232;input [7:0] in233;input [7:0] in234;input [7:0] in235;input [7:0] in236;input [7:0] in237;input [7:0] in238;input [7:0] in239;input [7:0] in240;input [7:0] in241;input [7:0] in242;input [7:0] in243;input [7:0] in244;input [7:0] in245;input [7:0] in246;input [7:0] in247;input [7:0] in248;input [7:0] in249;input [7:0] in250;input [7:0] in251;input [7:0] in252;input [7:0] in253;input [7:0] in254;input [7:0] in255;input [7:0] in256;input [7:0] in257;input [7:0] in258;input [7:0] in259;input [7:0] in260;input [7:0] in261;input [7:0] in262;input [7:0] in263;input [7:0] in264;input [7:0] in265;input [7:0] in266;input [7:0] in267;input [7:0] in268;input [7:0] in269;input [7:0] in270;input [7:0] in271;input [7:0] in272;input [7:0] in273;input [7:0] in274;input [7:0] in275;input [7:0] in276;input [7:0] in277;input [7:0] in278;input [7:0] in279;input [7:0] in280;input [7:0] in281;input [7:0] in282;input [7:0] in283;input [7:0] in284;input [7:0] in285;input [7:0] in286;input [7:0] in287;input [7:0] in288;input [7:0] in289;input [7:0] in290;input [7:0] in291;input [7:0] in292;input [7:0] in293;input [7:0] in294;input [7:0] in295;input [7:0] in296;input [7:0] in297;input [7:0] in298;input [7:0] in299;input [7:0] in300;input [7:0] in301;input [7:0] in302;input [7:0] in303;input [7:0] in304;input [7:0] in305;input [7:0] in306;input [7:0] in307;input [7:0] in308;input [7:0] in309;input [7:0] in310;input [7:0] in311;input [7:0] in312;input [7:0] in313;input [7:0] in314;input [7:0] in315;input [7:0] in316;input [7:0] in317;input [7:0] in318;input [7:0] in319;input [7:0] in320;input [7:0] in321;input [7:0] in322;input [7:0] in323;input [7:0] in324;input [7:0] in325;input [7:0] in326;input [7:0] in327;input [7:0] in328;input [7:0] in329;input [7:0] in330;input [7:0] in331;input [7:0] in332;input [7:0] in333;input [7:0] in334;input [7:0] in335;input [7:0] in336;input [7:0] in337;input [7:0] in338;input [7:0] in339;input [7:0] in340;input [7:0] in341;input [7:0] in342;input [7:0] in343;input [7:0] in344;input [7:0] in345;input [7:0] in346;input [7:0] in347;input [7:0] in348;input [7:0] in349;input [7:0] in350;input [7:0] in351;input [7:0] in352;input [7:0] in353;input [7:0] in354;input [7:0] in355;input [7:0] in356;input [7:0] in357;input [7:0] in358;input [7:0] in359;input [7:0] in360;input [7:0] in361;input [7:0] in362;input [7:0] in363;input [7:0] in364;input [7:0] in365;input [7:0] in366;input [7:0] in367;input [7:0] in368;input [7:0] in369;input [7:0] in370;input [7:0] in371;input [7:0] in372;input [7:0] in373;input [7:0] in374;input [7:0] in375;input [7:0] in376;input [7:0] in377;input [7:0] in378;input [7:0] in379;input [7:0] in380;input [7:0] in381;input [7:0] in382;input [7:0] in383;input [7:0] in384;input [7:0] in385;input [7:0] in386;input [7:0] in387;input [7:0] in388;input [7:0] in389;input [7:0] in390;input [7:0] in391;input [7:0] in392;input [7:0] in393;input [7:0] in394;input [7:0] in395;input [7:0] in396;input [7:0] in397;input [7:0] in398;input [7:0] in399;input [7:0] in400;input [7:0] in401;input [7:0] in402;input [7:0] in403;input [7:0] in404;input [7:0] in405;input [7:0] in406;input [7:0] in407;input [7:0] in408;input [7:0] in409;input [7:0] in410;input [7:0] in411;input [7:0] in412;input [7:0] in413;input [7:0] in414;input [7:0] in415;input [7:0] in416;input [7:0] in417;input [7:0] in418;input [7:0] in419;input [7:0] in420;input [7:0] in421;input [7:0] in422;input [7:0] in423;input [7:0] in424;input [7:0] in425;input [7:0] in426;input [7:0] in427;input [7:0] in428;input [7:0] in429;input [7:0] in430;input [7:0] in431;input [7:0] in432;input [7:0] in433;input [7:0] in434;input [7:0] in435;input [7:0] in436;input [7:0] in437;input [7:0] in438;input [7:0] in439;input [7:0] in440;input [7:0] in441;input [7:0] in442;input [7:0] in443;input [7:0] in444;input [7:0] in445;input [7:0] in446;input [7:0] in447;input [7:0] in448;input [7:0] in449;input [7:0] in450;input [7:0] in451;input [7:0] in452;input [7:0] in453;input [7:0] in454;input [7:0] in455;input [7:0] in456;input [7:0] in457;input [7:0] in458;input [7:0] in459;input [7:0] in460;input [7:0] in461;input [7:0] in462;input [7:0] in463;input [7:0] in464;input [7:0] in465;input [7:0] in466;input [7:0] in467;input [7:0] in468;input [7:0] in469;input [7:0] in470;input [7:0] in471;input [7:0] in472;input [7:0] in473;input [7:0] in474;input [7:0] in475;input [7:0] in476;input [7:0] in477;input [7:0] in478;input [7:0] in479;input [7:0] in480;input [7:0] in481;input [7:0] in482;input [7:0] in483;input [7:0] in484;input [7:0] in485;input [7:0] in486;input [7:0] in487;input [7:0] in488;input [7:0] in489;input [7:0] in490;input [7:0] in491;input [7:0] in492;input [7:0] in493;input [7:0] in494;input [7:0] in495;input [7:0] in496;input [7:0] in497;input [7:0] in498;input [7:0] in499;input [7:0] in500;input [7:0] in501;input [7:0] in502;input [7:0] in503;input [7:0] in504;input [7:0] in505;input [7:0] in506;input [7:0] in507;input [7:0] in508;input [7:0] in509;input [7:0] in510;input [7:0] in511;input [7:0] in512;input [7:0] in513;input [7:0] in514;input [7:0] in515;input [7:0] in516;input [7:0] in517;input [7:0] in518;input [7:0] in519;input [7:0] in520;input [7:0] in521;input [7:0] in522;input [7:0] in523;input [7:0] in524;input [7:0] in525;input [7:0] in526;input [7:0] in527;input [7:0] in528;input [7:0] in529;input [7:0] in530;input [7:0] in531;input [7:0] in532;input [7:0] in533;input [7:0] in534;input [7:0] in535;input [7:0] in536;input [7:0] in537;input [7:0] in538;input [7:0] in539;input [7:0] in540;input [7:0] in541;input [7:0] in542;input [7:0] in543;input [7:0] in544;input [7:0] in545;input [7:0] in546;input [7:0] in547;input [7:0] in548;input [7:0] in549;input [7:0] in550;input [7:0] in551;input [7:0] in552;input [7:0] in553;input [7:0] in554;input [7:0] in555;input [7:0] in556;input [7:0] in557;input [7:0] in558;input [7:0] in559;input [7:0] in560;input [7:0] in561;input [7:0] in562;input [7:0] in563;input [7:0] in564;input [7:0] in565;input [7:0] in566;input [7:0] in567;input [7:0] in568;input [7:0] in569;input [7:0] in570;input [7:0] in571;input [7:0] in572;input [7:0] in573;input [7:0] in574;input [7:0] in575;input [7:0] in576;input [7:0] in577;input [7:0] in578;input [7:0] in579;input [7:0] in580;input [7:0] in581;input [7:0] in582;input [7:0] in583;input [7:0] in584;input [7:0] in585;input [7:0] in586;input [7:0] in587;input [7:0] in588;input [7:0] in589;input [7:0] in590;input [7:0] in591;input [7:0] in592;input [7:0] in593;input [7:0] in594;input [7:0] in595;input [7:0] in596;input [7:0] in597;input [7:0] in598;input [7:0] in599;input [7:0] in600;input [7:0] in601;input [7:0] in602;input [7:0] in603;input [7:0] in604;input [7:0] in605;input [7:0] in606;input [7:0] in607;input [7:0] in608;input [7:0] in609;input [7:0] in610;input [7:0] in611;input [7:0] in612;input [7:0] in613;input [7:0] in614;input [7:0] in615;input [7:0] in616;input [7:0] in617;input [7:0] in618;input [7:0] in619;input [7:0] in620;input [7:0] in621;input [7:0] in622;input [7:0] in623;input [7:0] in624;input [7:0] in625;input [7:0] in626;input [7:0] in627;input [7:0] in628;input [7:0] in629;input [7:0] in630;input [7:0] in631;input [7:0] in632;input [7:0] in633;input [7:0] in634;input [7:0] in635;input [7:0] in636;input [7:0] in637;input [7:0] in638;input [7:0] in639;input [7:0] in640;input [7:0] in641;input [7:0] in642;input [7:0] in643;input [7:0] in644;input [7:0] in645;input [7:0] in646;input [7:0] in647;input [7:0] in648;input [7:0] in649;input [7:0] in650;input [7:0] in651;input [7:0] in652;input [7:0] in653;input [7:0] in654;input [7:0] in655;input [7:0] in656;input [7:0] in657;input [7:0] in658;input [7:0] in659;input [7:0] in660;input [7:0] in661;input [7:0] in662;input [7:0] in663;input [7:0] in664;input [7:0] in665;input [7:0] in666;input [7:0] in667;input [7:0] in668;input [7:0] in669;input [7:0] in670;input [7:0] in671;input [7:0] in672;input [7:0] in673;input [7:0] in674;input [7:0] in675;input [7:0] in676;input [7:0] in677;input [7:0] in678;input [7:0] in679;input [7:0] in680;input [7:0] in681;input [7:0] in682;input [7:0] in683;input [7:0] in684;input [7:0] in685;input [7:0] in686;input [7:0] in687;input [7:0] in688;input [7:0] in689;input [7:0] in690;input [7:0] in691;input [7:0] in692;input [7:0] in693;input [7:0] in694;input [7:0] in695;input [7:0] in696;input [7:0] in697;input [7:0] in698;input [7:0] in699;input [7:0] in700;input [7:0] in701;input [7:0] in702;input [7:0] in703;input [7:0] in704;input [7:0] in705;input [7:0] in706;input [7:0] in707;input [7:0] in708;input [7:0] in709;input [7:0] in710;input [7:0] in711;input [7:0] in712;input [7:0] in713;input [7:0] in714;input [7:0] in715;input [7:0] in716;input [7:0] in717;input [7:0] in718;input [7:0] in719;input [7:0] in720;input [7:0] in721;input [7:0] in722;input [7:0] in723;input [7:0] in724;input [7:0] in725;input [7:0] in726;input [7:0] in727;input [7:0] in728;input [7:0] in729;input [7:0] in730;input [7:0] in731;input [7:0] in732;input [7:0] in733;input [7:0] in734;input [7:0] in735;input [7:0] in736;input [7:0] in737;input [7:0] in738;input [7:0] in739;input [7:0] in740;input [7:0] in741;input [7:0] in742;input [7:0] in743;input [7:0] in744;input [7:0] in745;input [7:0] in746;input [7:0] in747;input [7:0] in748;input [7:0] in749;input [7:0] in750;input [7:0] in751;input [7:0] in752;input [7:0] in753;input [7:0] in754;input [7:0] in755;input [7:0] in756;input [7:0] in757;input [7:0] in758;input [7:0] in759;input [7:0] in760;input [7:0] in761;input [7:0] in762;input [7:0] in763;input [7:0] in764;input [7:0] in765;input [7:0] in766;input [7:0] in767;input [7:0] in768;input [7:0] in769;input [7:0] in770;input [7:0] in771;input [7:0] in772;input [7:0] in773;input [7:0] in774;input [7:0] in775;input [7:0] in776;input [7:0] in777;input [7:0] in778;input [7:0] in779;input [7:0] in780;input [7:0] in781;input [7:0] in782;input [7:0] in783;
input clk;input [7:0] bias;input start;output ready;output [7:0] out;

wire [7:0] con0;wire [7:0] con1;wire [7:0] con2;wire [7:0] con3;wire [7:0] con4;wire [7:0] con5;wire [7:0] con6;wire [7:0] con7;wire [7:0] con8;wire [7:0] con9;wire [7:0] con10;wire [7:0] con11;wire [7:0] con12;wire [7:0] con13;wire [7:0] con14;wire [7:0] con15;wire [7:0] con16;wire [7:0] con17;wire [7:0] con18;wire [7:0] con19;wire [7:0] con20;wire [7:0] con21;wire [7:0] con22;wire [7:0] con23;wire [7:0] con24;wire [7:0] con25;wire [7:0] con26;wire [7:0] con27;wire [7:0] con28;wire [7:0] con29;wire [7:0] con30;wire [7:0] con31;wire [7:0] con32;wire [7:0] con33;wire [7:0] con34;wire [7:0] con35;wire [7:0] con36;wire [7:0] con37;wire [7:0] con38;wire [7:0] con39;wire [7:0] con40;wire [7:0] con41;wire [7:0] con42;wire [7:0] con43;wire [7:0] con44;wire [7:0] con45;wire [7:0] con46;wire [7:0] con47;wire [7:0] con48;wire [7:0] con49;wire [7:0] con50;wire [7:0] con51;wire [7:0] con52;wire [7:0] con53;wire [7:0] con54;wire [7:0] con55;wire [7:0] con56;wire [7:0] con57;wire [7:0] con58;wire [7:0] con59;wire [7:0] con60;wire [7:0] con61;wire [7:0] con62;wire [7:0] con63;wire [7:0] con64;wire [7:0] con65;wire [7:0] con66;wire [7:0] con67;wire [7:0] con68;wire [7:0] con69;wire [7:0] con70;wire [7:0] con71;wire [7:0] con72;wire [7:0] con73;wire [7:0] con74;wire [7:0] con75;wire [7:0] con76;wire [7:0] con77;wire [7:0] con78;wire [7:0] con79;wire [7:0] con80;wire [7:0] con81;wire [7:0] con82;wire [7:0] con83;wire [7:0] con84;wire [7:0] con85;wire [7:0] con86;wire [7:0] con87;wire [7:0] con88;wire [7:0] con89;wire [7:0] con90;wire [7:0] con91;wire [7:0] con92;wire [7:0] con93;wire [7:0] con94;wire [7:0] con95;wire [7:0] con96;wire [7:0] con97;wire [7:0] con98;wire [7:0] con99;wire [7:0] con100;wire [7:0] con101;wire [7:0] con102;wire [7:0] con103;wire [7:0] con104;wire [7:0] con105;wire [7:0] con106;wire [7:0] con107;wire [7:0] con108;wire [7:0] con109;wire [7:0] con110;wire [7:0] con111;wire [7:0] con112;wire [7:0] con113;wire [7:0] con114;wire [7:0] con115;wire [7:0] con116;wire [7:0] con117;wire [7:0] con118;wire [7:0] con119;wire [7:0] con120;wire [7:0] con121;wire [7:0] con122;wire [7:0] con123;wire [7:0] con124;wire [7:0] con125;wire [7:0] con126;wire [7:0] con127;wire [7:0] con128;wire [7:0] con129;wire [7:0] con130;wire [7:0] con131;wire [7:0] con132;wire [7:0] con133;wire [7:0] con134;wire [7:0] con135;wire [7:0] con136;wire [7:0] con137;wire [7:0] con138;wire [7:0] con139;wire [7:0] con140;wire [7:0] con141;wire [7:0] con142;wire [7:0] con143;wire [7:0] con144;wire [7:0] con145;wire [7:0] con146;wire [7:0] con147;wire [7:0] con148;wire [7:0] con149;wire [7:0] con150;wire [7:0] con151;wire [7:0] con152;wire [7:0] con153;wire [7:0] con154;wire [7:0] con155;wire [7:0] con156;wire [7:0] con157;wire [7:0] con158;wire [7:0] con159;wire [7:0] con160;wire [7:0] con161;wire [7:0] con162;wire [7:0] con163;wire [7:0] con164;wire [7:0] con165;wire [7:0] con166;wire [7:0] con167;wire [7:0] con168;wire [7:0] con169;wire [7:0] con170;wire [7:0] con171;wire [7:0] con172;wire [7:0] con173;wire [7:0] con174;wire [7:0] con175;wire [7:0] con176;wire [7:0] con177;wire [7:0] con178;wire [7:0] con179;wire [7:0] con180;wire [7:0] con181;wire [7:0] con182;wire [7:0] con183;wire [7:0] con184;wire [7:0] con185;wire [7:0] con186;wire [7:0] con187;wire [7:0] con188;wire [7:0] con189;wire [7:0] con190;wire [7:0] con191;wire [7:0] con192;wire [7:0] con193;wire [7:0] con194;wire [7:0] con195;wire [7:0] con196;wire [7:0] con197;wire [7:0] con198;wire [7:0] con199;wire [7:0] con200;wire [7:0] con201;wire [7:0] con202;wire [7:0] con203;wire [7:0] con204;wire [7:0] con205;wire [7:0] con206;wire [7:0] con207;wire [7:0] con208;wire [7:0] con209;wire [7:0] con210;wire [7:0] con211;wire [7:0] con212;wire [7:0] con213;wire [7:0] con214;wire [7:0] con215;wire [7:0] con216;wire [7:0] con217;wire [7:0] con218;wire [7:0] con219;wire [7:0] con220;wire [7:0] con221;wire [7:0] con222;wire [7:0] con223;wire [7:0] con224;wire [7:0] con225;wire [7:0] con226;wire [7:0] con227;wire [7:0] con228;wire [7:0] con229;wire [7:0] con230;wire [7:0] con231;wire [7:0] con232;wire [7:0] con233;wire [7:0] con234;wire [7:0] con235;wire [7:0] con236;wire [7:0] con237;wire [7:0] con238;wire [7:0] con239;wire [7:0] con240;wire [7:0] con241;wire [7:0] con242;wire [7:0] con243;wire [7:0] con244;wire [7:0] con245;wire [7:0] con246;wire [7:0] con247;wire [7:0] con248;wire [7:0] con249;wire [7:0] con250;wire [7:0] con251;wire [7:0] con252;wire [7:0] con253;wire [7:0] con254;wire [7:0] con255;wire [7:0] con256;wire [7:0] con257;wire [7:0] con258;wire [7:0] con259;wire [7:0] con260;wire [7:0] con261;wire [7:0] con262;wire [7:0] con263;wire [7:0] con264;wire [7:0] con265;wire [7:0] con266;wire [7:0] con267;wire [7:0] con268;wire [7:0] con269;wire [7:0] con270;wire [7:0] con271;wire [7:0] con272;wire [7:0] con273;wire [7:0] con274;wire [7:0] con275;wire [7:0] con276;wire [7:0] con277;wire [7:0] con278;wire [7:0] con279;wire [7:0] con280;wire [7:0] con281;wire [7:0] con282;wire [7:0] con283;wire [7:0] con284;wire [7:0] con285;wire [7:0] con286;wire [7:0] con287;wire [7:0] con288;wire [7:0] con289;wire [7:0] con290;wire [7:0] con291;wire [7:0] con292;wire [7:0] con293;wire [7:0] con294;wire [7:0] con295;wire [7:0] con296;wire [7:0] con297;wire [7:0] con298;wire [7:0] con299;wire [7:0] con300;wire [7:0] con301;wire [7:0] con302;wire [7:0] con303;wire [7:0] con304;wire [7:0] con305;wire [7:0] con306;wire [7:0] con307;wire [7:0] con308;wire [7:0] con309;wire [7:0] con310;wire [7:0] con311;wire [7:0] con312;wire [7:0] con313;wire [7:0] con314;wire [7:0] con315;wire [7:0] con316;wire [7:0] con317;wire [7:0] con318;wire [7:0] con319;wire [7:0] con320;wire [7:0] con321;wire [7:0] con322;wire [7:0] con323;wire [7:0] con324;wire [7:0] con325;wire [7:0] con326;wire [7:0] con327;wire [7:0] con328;wire [7:0] con329;wire [7:0] con330;wire [7:0] con331;wire [7:0] con332;wire [7:0] con333;wire [7:0] con334;wire [7:0] con335;wire [7:0] con336;wire [7:0] con337;wire [7:0] con338;wire [7:0] con339;wire [7:0] con340;wire [7:0] con341;wire [7:0] con342;wire [7:0] con343;wire [7:0] con344;wire [7:0] con345;wire [7:0] con346;wire [7:0] con347;wire [7:0] con348;wire [7:0] con349;wire [7:0] con350;wire [7:0] con351;wire [7:0] con352;wire [7:0] con353;wire [7:0] con354;wire [7:0] con355;wire [7:0] con356;wire [7:0] con357;wire [7:0] con358;wire [7:0] con359;wire [7:0] con360;wire [7:0] con361;wire [7:0] con362;wire [7:0] con363;wire [7:0] con364;wire [7:0] con365;wire [7:0] con366;wire [7:0] con367;wire [7:0] con368;wire [7:0] con369;wire [7:0] con370;wire [7:0] con371;wire [7:0] con372;wire [7:0] con373;wire [7:0] con374;wire [7:0] con375;wire [7:0] con376;wire [7:0] con377;wire [7:0] con378;wire [7:0] con379;wire [7:0] con380;wire [7:0] con381;wire [7:0] con382;wire [7:0] con383;wire [7:0] con384;wire [7:0] con385;wire [7:0] con386;wire [7:0] con387;wire [7:0] con388;wire [7:0] con389;wire [7:0] con390;wire [7:0] con391;wire [7:0] con392;wire [7:0] con393;wire [7:0] con394;wire [7:0] con395;wire [7:0] con396;wire [7:0] con397;wire [7:0] con398;wire [7:0] con399;wire [7:0] con400;wire [7:0] con401;wire [7:0] con402;wire [7:0] con403;wire [7:0] con404;wire [7:0] con405;wire [7:0] con406;wire [7:0] con407;wire [7:0] con408;wire [7:0] con409;wire [7:0] con410;wire [7:0] con411;wire [7:0] con412;wire [7:0] con413;wire [7:0] con414;wire [7:0] con415;wire [7:0] con416;wire [7:0] con417;wire [7:0] con418;wire [7:0] con419;wire [7:0] con420;wire [7:0] con421;wire [7:0] con422;wire [7:0] con423;wire [7:0] con424;wire [7:0] con425;wire [7:0] con426;wire [7:0] con427;wire [7:0] con428;wire [7:0] con429;wire [7:0] con430;wire [7:0] con431;wire [7:0] con432;wire [7:0] con433;wire [7:0] con434;wire [7:0] con435;wire [7:0] con436;wire [7:0] con437;wire [7:0] con438;wire [7:0] con439;wire [7:0] con440;wire [7:0] con441;wire [7:0] con442;wire [7:0] con443;wire [7:0] con444;wire [7:0] con445;wire [7:0] con446;wire [7:0] con447;wire [7:0] con448;wire [7:0] con449;wire [7:0] con450;wire [7:0] con451;wire [7:0] con452;wire [7:0] con453;wire [7:0] con454;wire [7:0] con455;wire [7:0] con456;wire [7:0] con457;wire [7:0] con458;wire [7:0] con459;wire [7:0] con460;wire [7:0] con461;wire [7:0] con462;wire [7:0] con463;wire [7:0] con464;wire [7:0] con465;wire [7:0] con466;wire [7:0] con467;wire [7:0] con468;wire [7:0] con469;wire [7:0] con470;wire [7:0] con471;wire [7:0] con472;wire [7:0] con473;wire [7:0] con474;wire [7:0] con475;wire [7:0] con476;wire [7:0] con477;wire [7:0] con478;wire [7:0] con479;wire [7:0] con480;wire [7:0] con481;wire [7:0] con482;wire [7:0] con483;wire [7:0] con484;wire [7:0] con485;wire [7:0] con486;wire [7:0] con487;wire [7:0] con488;wire [7:0] con489;wire [7:0] con490;wire [7:0] con491;wire [7:0] con492;wire [7:0] con493;wire [7:0] con494;wire [7:0] con495;wire [7:0] con496;wire [7:0] con497;wire [7:0] con498;wire [7:0] con499;wire [7:0] con500;wire [7:0] con501;wire [7:0] con502;wire [7:0] con503;wire [7:0] con504;wire [7:0] con505;wire [7:0] con506;wire [7:0] con507;wire [7:0] con508;wire [7:0] con509;wire [7:0] con510;wire [7:0] con511;wire [7:0] con512;wire [7:0] con513;wire [7:0] con514;wire [7:0] con515;wire [7:0] con516;wire [7:0] con517;wire [7:0] con518;wire [7:0] con519;wire [7:0] con520;wire [7:0] con521;wire [7:0] con522;wire [7:0] con523;wire [7:0] con524;wire [7:0] con525;wire [7:0] con526;wire [7:0] con527;wire [7:0] con528;wire [7:0] con529;wire [7:0] con530;wire [7:0] con531;wire [7:0] con532;wire [7:0] con533;wire [7:0] con534;wire [7:0] con535;wire [7:0] con536;wire [7:0] con537;wire [7:0] con538;wire [7:0] con539;wire [7:0] con540;wire [7:0] con541;wire [7:0] con542;wire [7:0] con543;wire [7:0] con544;wire [7:0] con545;wire [7:0] con546;wire [7:0] con547;wire [7:0] con548;wire [7:0] con549;wire [7:0] con550;wire [7:0] con551;wire [7:0] con552;wire [7:0] con553;wire [7:0] con554;wire [7:0] con555;wire [7:0] con556;wire [7:0] con557;wire [7:0] con558;wire [7:0] con559;wire [7:0] con560;wire [7:0] con561;wire [7:0] con562;wire [7:0] con563;wire [7:0] con564;wire [7:0] con565;wire [7:0] con566;wire [7:0] con567;wire [7:0] con568;wire [7:0] con569;wire [7:0] con570;wire [7:0] con571;wire [7:0] con572;wire [7:0] con573;wire [7:0] con574;wire [7:0] con575;
wire readycon;wire readypool; 

ConvLayer conl1(.weight0(weight1l0),.weight1(weight1l1),.weight2(weight1l2),.weight3(weight1l3),.weight4(weight1l4),.weight5(weight1l5),.weight6(weight1l6),.weight7(weight1l7),.weight8(weight1l8),.weight9(weight1l9),.weight10(weight1l10),.weight11(weight1l11),.weight12(weight1l12),.weight13(weight1l13),.weight14(weight1l14),.weight15(weight1l15),.weight16(weight1l16),.weight17(weight1l17),.weight18(weight1l18),.weight19(weight1l19),.weight20(weight1l20),.weight21(weight1l21),.weight22(weight1l22),.weight23(weight1l23),.weight24(weight1l24),
.in0(in0),.in1(in1),.in2(in2),.in3(in3),.in4(in4),.in5(in5),.in6(in6),.in7(in7),.in8(in8),.in9(in9),.in10(in10),.in11(in11),.in12(in12),.in13(in13),.in14(in14),.in15(in15),.in16(in16),.in17(in17),.in18(in18),.in19(in19),.in20(in20),.in21(in21),.in22(in22),.in23(in23),.in24(in24),.in25(in25),.in26(in26),.in27(in27),.in28(in28),.in29(in29),.in30(in30),.in31(in31),.in32(in32),.in33(in33),.in34(in34),.in35(in35),.in36(in36),.in37(in37),.in38(in38),.in39(in39),.in40(in40),.in41(in41),.in42(in42),.in43(in43),.in44(in44),.in45(in45),.in46(in46),.in47(in47),.in48(in48),.in49(in49),.in50(in50),.in51(in51),.in52(in52),.in53(in53),.in54(in54),.in55(in55),.in56(in56),.in57(in57),.in58(in58),.in59(in59),.in60(in60),.in61(in61),.in62(in62),.in63(in63),.in64(in64),.in65(in65),.in66(in66),.in67(in67),.in68(in68),.in69(in69),.in70(in70),.in71(in71),.in72(in72),.in73(in73),.in74(in74),.in75(in75),.in76(in76),.in77(in77),.in78(in78),.in79(in79),.in80(in80),.in81(in81),.in82(in82),.in83(in83),.in84(in84),.in85(in85),.in86(in86),.in87(in87),.in88(in88),.in89(in89),.in90(in90),.in91(in91),.in92(in92),.in93(in93),.in94(in94),.in95(in95),.in96(in96),.in97(in97),.in98(in98),.in99(in99),.in100(in100),.in101(in101),.in102(in102),.in103(in103),.in104(in104),.in105(in105),.in106(in106),.in107(in107),.in108(in108),.in109(in109),.in110(in110),.in111(in111),.in112(in112),.in113(in113),.in114(in114),.in115(in115),.in116(in116),.in117(in117),.in118(in118),.in119(in119),.in120(in120),.in121(in121),.in122(in122),.in123(in123),.in124(in124),.in125(in125),.in126(in126),.in127(in127),.in128(in128),.in129(in129),.in130(in130),.in131(in131),.in132(in132),.in133(in133),.in134(in134),.in135(in135),.in136(in136),.in137(in137),.in138(in138),.in139(in139),.in140(in140),.in141(in141),.in142(in142),.in143(in143),.in144(in144),.in145(in145),.in146(in146),.in147(in147),.in148(in148),.in149(in149),.in150(in150),.in151(in151),.in152(in152),.in153(in153),.in154(in154),.in155(in155),.in156(in156),.in157(in157),.in158(in158),.in159(in159),.in160(in160),.in161(in161),.in162(in162),.in163(in163),.in164(in164),.in165(in165),.in166(in166),.in167(in167),.in168(in168),.in169(in169),.in170(in170),.in171(in171),.in172(in172),.in173(in173),.in174(in174),.in175(in175),.in176(in176),.in177(in177),.in178(in178),.in179(in179),.in180(in180),.in181(in181),.in182(in182),.in183(in183),.in184(in184),.in185(in185),.in186(in186),.in187(in187),.in188(in188),.in189(in189),.in190(in190),.in191(in191),.in192(in192),.in193(in193),.in194(in194),.in195(in195),.in196(in196),.in197(in197),.in198(in198),.in199(in199),.in200(in200),.in201(in201),.in202(in202),.in203(in203),.in204(in204),.in205(in205),.in206(in206),.in207(in207),.in208(in208),.in209(in209),.in210(in210),.in211(in211),.in212(in212),.in213(in213),.in214(in214),.in215(in215),.in216(in216),.in217(in217),.in218(in218),.in219(in219),.in220(in220),.in221(in221),.in222(in222),.in223(in223),.in224(in224),.in225(in225),.in226(in226),.in227(in227),.in228(in228),.in229(in229),.in230(in230),.in231(in231),.in232(in232),.in233(in233),.in234(in234),.in235(in235),.in236(in236),.in237(in237),.in238(in238),.in239(in239),.in240(in240),.in241(in241),.in242(in242),.in243(in243),.in244(in244),.in245(in245),.in246(in246),.in247(in247),.in248(in248),.in249(in249),.in250(in250),.in251(in251),.in252(in252),.in253(in253),.in254(in254),.in255(in255),.in256(in256),.in257(in257),.in258(in258),.in259(in259),.in260(in260),.in261(in261),.in262(in262),.in263(in263),.in264(in264),.in265(in265),.in266(in266),.in267(in267),.in268(in268),.in269(in269),.in270(in270),.in271(in271),.in272(in272),.in273(in273),.in274(in274),.in275(in275),.in276(in276),.in277(in277),.in278(in278),.in279(in279),.in280(in280),.in281(in281),.in282(in282),.in283(in283),.in284(in284),.in285(in285),.in286(in286),.in287(in287),.in288(in288),.in289(in289),.in290(in290),.in291(in291),.in292(in292),.in293(in293),.in294(in294),.in295(in295),.in296(in296),.in297(in297),.in298(in298),.in299(in299),.in300(in300),.in301(in301),.in302(in302),.in303(in303),.in304(in304),.in305(in305),.in306(in306),.in307(in307),.in308(in308),.in309(in309),.in310(in310),.in311(in311),.in312(in312),.in313(in313),.in314(in314),.in315(in315),.in316(in316),.in317(in317),.in318(in318),.in319(in319),.in320(in320),.in321(in321),.in322(in322),.in323(in323),.in324(in324),.in325(in325),.in326(in326),.in327(in327),.in328(in328),.in329(in329),.in330(in330),.in331(in331),.in332(in332),.in333(in333),.in334(in334),.in335(in335),.in336(in336),.in337(in337),.in338(in338),.in339(in339),.in340(in340),.in341(in341),.in342(in342),.in343(in343),.in344(in344),.in345(in345),.in346(in346),.in347(in347),.in348(in348),.in349(in349),.in350(in350),.in351(in351),.in352(in352),.in353(in353),.in354(in354),.in355(in355),.in356(in356),.in357(in357),.in358(in358),.in359(in359),.in360(in360),.in361(in361),.in362(in362),.in363(in363),.in364(in364),.in365(in365),.in366(in366),.in367(in367),.in368(in368),.in369(in369),.in370(in370),.in371(in371),.in372(in372),.in373(in373),.in374(in374),.in375(in375),.in376(in376),.in377(in377),.in378(in378),.in379(in379),.in380(in380),.in381(in381),.in382(in382),.in383(in383),.in384(in384),.in385(in385),.in386(in386),.in387(in387),.in388(in388),.in389(in389),.in390(in390),.in391(in391),.in392(in392),.in393(in393),.in394(in394),.in395(in395),.in396(in396),.in397(in397),.in398(in398),.in399(in399),.in400(in400),.in401(in401),.in402(in402),.in403(in403),.in404(in404),.in405(in405),.in406(in406),.in407(in407),.in408(in408),.in409(in409),.in410(in410),.in411(in411),.in412(in412),.in413(in413),.in414(in414),.in415(in415),.in416(in416),.in417(in417),.in418(in418),.in419(in419),.in420(in420),.in421(in421),.in422(in422),.in423(in423),.in424(in424),.in425(in425),.in426(in426),.in427(in427),.in428(in428),.in429(in429),.in430(in430),.in431(in431),.in432(in432),.in433(in433),.in434(in434),.in435(in435),.in436(in436),.in437(in437),.in438(in438),.in439(in439),.in440(in440),.in441(in441),.in442(in442),.in443(in443),.in444(in444),.in445(in445),.in446(in446),.in447(in447),.in448(in448),.in449(in449),.in450(in450),.in451(in451),.in452(in452),.in453(in453),.in454(in454),.in455(in455),.in456(in456),.in457(in457),.in458(in458),.in459(in459),.in460(in460),.in461(in461),.in462(in462),.in463(in463),.in464(in464),.in465(in465),.in466(in466),.in467(in467),.in468(in468),.in469(in469),.in470(in470),.in471(in471),.in472(in472),.in473(in473),.in474(in474),.in475(in475),.in476(in476),.in477(in477),.in478(in478),.in479(in479),.in480(in480),.in481(in481),.in482(in482),.in483(in483),.in484(in484),.in485(in485),.in486(in486),.in487(in487),.in488(in488),.in489(in489),.in490(in490),.in491(in491),.in492(in492),.in493(in493),.in494(in494),.in495(in495),.in496(in496),.in497(in497),.in498(in498),.in499(in499),.in500(in500),.in501(in501),.in502(in502),.in503(in503),.in504(in504),.in505(in505),.in506(in506),.in507(in507),.in508(in508),.in509(in509),.in510(in510),.in511(in511),.in512(in512),.in513(in513),.in514(in514),.in515(in515),.in516(in516),.in517(in517),.in518(in518),.in519(in519),.in520(in520),.in521(in521),.in522(in522),.in523(in523),.in524(in524),.in525(in525),.in526(in526),.in527(in527),.in528(in528),.in529(in529),.in530(in530),.in531(in531),.in532(in532),.in533(in533),.in534(in534),.in535(in535),.in536(in536),.in537(in537),.in538(in538),.in539(in539),.in540(in540),.in541(in541),.in542(in542),.in543(in543),.in544(in544),.in545(in545),.in546(in546),.in547(in547),.in548(in548),.in549(in549),.in550(in550),.in551(in551),.in552(in552),.in553(in553),.in554(in554),.in555(in555),.in556(in556),.in557(in557),.in558(in558),.in559(in559),.in560(in560),.in561(in561),.in562(in562),.in563(in563),.in564(in564),.in565(in565),.in566(in566),.in567(in567),.in568(in568),.in569(in569),.in570(in570),.in571(in571),.in572(in572),.in573(in573),.in574(in574),.in575(in575),.in576(in576),.in577(in577),.in578(in578),.in579(in579),.in580(in580),.in581(in581),.in582(in582),.in583(in583),.in584(in584),.in585(in585),.in586(in586),.in587(in587),.in588(in588),.in589(in589),.in590(in590),.in591(in591),.in592(in592),.in593(in593),.in594(in594),.in595(in595),.in596(in596),.in597(in597),.in598(in598),.in599(in599),.in600(in600),.in601(in601),.in602(in602),.in603(in603),.in604(in604),.in605(in605),.in606(in606),.in607(in607),.in608(in608),.in609(in609),.in610(in610),.in611(in611),.in612(in612),.in613(in613),.in614(in614),.in615(in615),.in616(in616),.in617(in617),.in618(in618),.in619(in619),.in620(in620),.in621(in621),.in622(in622),.in623(in623),.in624(in624),.in625(in625),.in626(in626),.in627(in627),.in628(in628),.in629(in629),.in630(in630),.in631(in631),.in632(in632),.in633(in633),.in634(in634),.in635(in635),.in636(in636),.in637(in637),.in638(in638),.in639(in639),.in640(in640),.in641(in641),.in642(in642),.in643(in643),.in644(in644),.in645(in645),.in646(in646),.in647(in647),.in648(in648),.in649(in649),.in650(in650),.in651(in651),.in652(in652),.in653(in653),.in654(in654),.in655(in655),.in656(in656),.in657(in657),.in658(in658),.in659(in659),.in660(in660),.in661(in661),.in662(in662),.in663(in663),.in664(in664),.in665(in665),.in666(in666),.in667(in667),.in668(in668),.in669(in669),.in670(in670),.in671(in671),.in672(in672),.in673(in673),.in674(in674),.in675(in675),.in676(in676),.in677(in677),.in678(in678),.in679(in679),.in680(in680),.in681(in681),.in682(in682),.in683(in683),.in684(in684),.in685(in685),.in686(in686),.in687(in687),.in688(in688),.in689(in689),.in690(in690),.in691(in691),.in692(in692),.in693(in693),.in694(in694),.in695(in695),.in696(in696),.in697(in697),.in698(in698),.in699(in699),.in700(in700),.in701(in701),.in702(in702),.in703(in703),.in704(in704),.in705(in705),.in706(in706),.in707(in707),.in708(in708),.in709(in709),.in710(in710),.in711(in711),.in712(in712),.in713(in713),.in714(in714),.in715(in715),.in716(in716),.in717(in717),.in718(in718),.in719(in719),.in720(in720),.in721(in721),.in722(in722),.in723(in723),.in724(in724),.in725(in725),.in726(in726),.in727(in727),.in728(in728),.in729(in729),.in730(in730),.in731(in731),.in732(in732),.in733(in733),.in734(in734),.in735(in735),.in736(in736),.in737(in737),.in738(in738),.in739(in739),.in740(in740),.in741(in741),.in742(in742),.in743(in743),.in744(in744),.in745(in745),.in746(in746),.in747(in747),.in748(in748),.in749(in749),.in750(in750),.in751(in751),.in752(in752),.in753(in753),.in754(in754),.in755(in755),.in756(in756),.in757(in757),.in758(in758),.in759(in759),.in760(in760),.in761(in761),.in762(in762),.in763(in763),.in764(in764),.in765(in765),.in766(in766),.in767(in767),.in768(in768),.in769(in769),.in770(in770),.in771(in771),.in772(in772),.in773(in773),.in774(in774),.in775(in775),.in776(in776),.in777(in777),.in778(in778),.in779(in779),.in780(in780),.in781(in781),.in782(in782),.in783(in783),
.conv0(con0),.conv1(con1),.conv2(con2),.conv3(con3),.conv4(con4),.conv5(con5),.conv6(con6),.conv7(con7),.conv8(con8),.conv9(con9),.conv10(con10),.conv11(con11),.conv12(con12),.conv13(con13),.conv14(con14),.conv15(con15),.conv16(con16),.conv17(con17),.conv18(con18),.conv19(con19),.conv20(con20),.conv21(con21),.conv22(con22),.conv23(con23),.conv24(con24),.conv25(con25),.conv26(con26),.conv27(con27),.conv28(con28),.conv29(con29),.conv30(con30),.conv31(con31),.conv32(con32),.conv33(con33),.conv34(con34),.conv35(con35),.conv36(con36),.conv37(con37),.conv38(con38),.conv39(con39),.conv40(con40),.conv41(con41),.conv42(con42),.conv43(con43),.conv44(con44),.conv45(con45),.conv46(con46),.conv47(con47),.conv48(con48),.conv49(con49),.conv50(con50),.conv51(con51),.conv52(con52),.conv53(con53),.conv54(con54),.conv55(con55),.conv56(con56),.conv57(con57),.conv58(con58),.conv59(con59),.conv60(con60),.conv61(con61),.conv62(con62),.conv63(con63),.conv64(con64),.conv65(con65),.conv66(con66),.conv67(con67),.conv68(con68),.conv69(con69),.conv70(con70),.conv71(con71),.conv72(con72),.conv73(con73),.conv74(con74),.conv75(con75),.conv76(con76),.conv77(con77),.conv78(con78),.conv79(con79),.conv80(con80),.conv81(con81),.conv82(con82),.conv83(con83),.conv84(con84),.conv85(con85),.conv86(con86),.conv87(con87),.conv88(con88),.conv89(con89),.conv90(con90),.conv91(con91),.conv92(con92),.conv93(con93),.conv94(con94),.conv95(con95),.conv96(con96),.conv97(con97),.conv98(con98),.conv99(con99),.conv100(con100),.conv101(con101),.conv102(con102),.conv103(con103),.conv104(con104),.conv105(con105),.conv106(con106),.conv107(con107),.conv108(con108),.conv109(con109),.conv110(con110),.conv111(con111),.conv112(con112),.conv113(con113),.conv114(con114),.conv115(con115),.conv116(con116),.conv117(con117),.conv118(con118),.conv119(con119),.conv120(con120),.conv121(con121),.conv122(con122),.conv123(con123),.conv124(con124),.conv125(con125),.conv126(con126),.conv127(con127),.conv128(con128),.conv129(con129),.conv130(con130),.conv131(con131),.conv132(con132),.conv133(con133),.conv134(con134),.conv135(con135),.conv136(con136),.conv137(con137),.conv138(con138),.conv139(con139),.conv140(con140),.conv141(con141),.conv142(con142),.conv143(con143),.conv144(con144),.conv145(con145),.conv146(con146),.conv147(con147),.conv148(con148),.conv149(con149),.conv150(con150),.conv151(con151),.conv152(con152),.conv153(con153),.conv154(con154),.conv155(con155),.conv156(con156),.conv157(con157),.conv158(con158),.conv159(con159),.conv160(con160),.conv161(con161),.conv162(con162),.conv163(con163),.conv164(con164),.conv165(con165),.conv166(con166),.conv167(con167),.conv168(con168),.conv169(con169),.conv170(con170),.conv171(con171),.conv172(con172),.conv173(con173),.conv174(con174),.conv175(con175),.conv176(con176),.conv177(con177),.conv178(con178),.conv179(con179),.conv180(con180),.conv181(con181),.conv182(con182),.conv183(con183),.conv184(con184),.conv185(con185),.conv186(con186),.conv187(con187),.conv188(con188),.conv189(con189),.conv190(con190),.conv191(con191),.conv192(con192),.conv193(con193),.conv194(con194),.conv195(con195),.conv196(con196),.conv197(con197),.conv198(con198),.conv199(con199),.conv200(con200),.conv201(con201),.conv202(con202),.conv203(con203),.conv204(con204),.conv205(con205),.conv206(con206),.conv207(con207),.conv208(con208),.conv209(con209),.conv210(con210),.conv211(con211),.conv212(con212),.conv213(con213),.conv214(con214),.conv215(con215),.conv216(con216),.conv217(con217),.conv218(con218),.conv219(con219),.conv220(con220),.conv221(con221),.conv222(con222),.conv223(con223),.conv224(con224),.conv225(con225),.conv226(con226),.conv227(con227),.conv228(con228),.conv229(con229),.conv230(con230),.conv231(con231),.conv232(con232),.conv233(con233),.conv234(con234),.conv235(con235),.conv236(con236),.conv237(con237),.conv238(con238),.conv239(con239),.conv240(con240),.conv241(con241),.conv242(con242),.conv243(con243),.conv244(con244),.conv245(con245),.conv246(con246),.conv247(con247),.conv248(con248),.conv249(con249),.conv250(con250),.conv251(con251),.conv252(con252),.conv253(con253),.conv254(con254),.conv255(con255),.conv256(con256),.conv257(con257),.conv258(con258),.conv259(con259),.conv260(con260),.conv261(con261),.conv262(con262),.conv263(con263),.conv264(con264),.conv265(con265),.conv266(con266),.conv267(con267),.conv268(con268),.conv269(con269),.conv270(con270),.conv271(con271),.conv272(con272),.conv273(con273),.conv274(con274),.conv275(con275),.conv276(con276),.conv277(con277),.conv278(con278),.conv279(con279),.conv280(con280),.conv281(con281),.conv282(con282),.conv283(con283),.conv284(con284),.conv285(con285),.conv286(con286),.conv287(con287),.conv288(con288),.conv289(con289),.conv290(con290),.conv291(con291),.conv292(con292),.conv293(con293),.conv294(con294),.conv295(con295),.conv296(con296),.conv297(con297),.conv298(con298),.conv299(con299),.conv300(con300),.conv301(con301),.conv302(con302),.conv303(con303),.conv304(con304),.conv305(con305),.conv306(con306),.conv307(con307),.conv308(con308),.conv309(con309),.conv310(con310),.conv311(con311),.conv312(con312),.conv313(con313),.conv314(con314),.conv315(con315),.conv316(con316),.conv317(con317),.conv318(con318),.conv319(con319),.conv320(con320),.conv321(con321),.conv322(con322),.conv323(con323),.conv324(con324),.conv325(con325),.conv326(con326),.conv327(con327),.conv328(con328),.conv329(con329),.conv330(con330),.conv331(con331),.conv332(con332),.conv333(con333),.conv334(con334),.conv335(con335),.conv336(con336),.conv337(con337),.conv338(con338),.conv339(con339),.conv340(con340),.conv341(con341),.conv342(con342),.conv343(con343),.conv344(con344),.conv345(con345),.conv346(con346),.conv347(con347),.conv348(con348),.conv349(con349),.conv350(con350),.conv351(con351),.conv352(con352),.conv353(con353),.conv354(con354),.conv355(con355),.conv356(con356),.conv357(con357),.conv358(con358),.conv359(con359),.conv360(con360),.conv361(con361),.conv362(con362),.conv363(con363),.conv364(con364),.conv365(con365),.conv366(con366),.conv367(con367),.conv368(con368),.conv369(con369),.conv370(con370),.conv371(con371),.conv372(con372),.conv373(con373),.conv374(con374),.conv375(con375),.conv376(con376),.conv377(con377),.conv378(con378),.conv379(con379),.conv380(con380),.conv381(con381),.conv382(con382),.conv383(con383),.conv384(con384),.conv385(con385),.conv386(con386),.conv387(con387),.conv388(con388),.conv389(con389),.conv390(con390),.conv391(con391),.conv392(con392),.conv393(con393),.conv394(con394),.conv395(con395),.conv396(con396),.conv397(con397),.conv398(con398),.conv399(con399),.conv400(con400),.conv401(con401),.conv402(con402),.conv403(con403),.conv404(con404),.conv405(con405),.conv406(con406),.conv407(con407),.conv408(con408),.conv409(con409),.conv410(con410),.conv411(con411),.conv412(con412),.conv413(con413),.conv414(con414),.conv415(con415),.conv416(con416),.conv417(con417),.conv418(con418),.conv419(con419),.conv420(con420),.conv421(con421),.conv422(con422),.conv423(con423),.conv424(con424),.conv425(con425),.conv426(con426),.conv427(con427),.conv428(con428),.conv429(con429),.conv430(con430),.conv431(con431),.conv432(con432),.conv433(con433),.conv434(con434),.conv435(con435),.conv436(con436),.conv437(con437),.conv438(con438),.conv439(con439),.conv440(con440),.conv441(con441),.conv442(con442),.conv443(con443),.conv444(con444),.conv445(con445),.conv446(con446),.conv447(con447),.conv448(con448),.conv449(con449),.conv450(con450),.conv451(con451),.conv452(con452),.conv453(con453),.conv454(con454),.conv455(con455),.conv456(con456),.conv457(con457),.conv458(con458),.conv459(con459),.conv460(con460),.conv461(con461),.conv462(con462),.conv463(con463),.conv464(con464),.conv465(con465),.conv466(con466),.conv467(con467),.conv468(con468),.conv469(con469),.conv470(con470),.conv471(con471),.conv472(con472),.conv473(con473),.conv474(con474),.conv475(con475),.conv476(con476),.conv477(con477),.conv478(con478),.conv479(con479),.conv480(con480),.conv481(con481),.conv482(con482),.conv483(con483),.conv484(con484),.conv485(con485),.conv486(con486),.conv487(con487),.conv488(con488),.conv489(con489),.conv490(con490),.conv491(con491),.conv492(con492),.conv493(con493),.conv494(con494),.conv495(con495),.conv496(con496),.conv497(con497),.conv498(con498),.conv499(con499),.conv500(con500),.conv501(con501),.conv502(con502),.conv503(con503),.conv504(con504),.conv505(con505),.conv506(con506),.conv507(con507),.conv508(con508),.conv509(con509),.conv510(con510),.conv511(con511),.conv512(con512),.conv513(con513),.conv514(con514),.conv515(con515),.conv516(con516),.conv517(con517),.conv518(con518),.conv519(con519),.conv520(con520),.conv521(con521),.conv522(con522),.conv523(con523),.conv524(con524),.conv525(con525),.conv526(con526),.conv527(con527),.conv528(con528),.conv529(con529),.conv530(con530),.conv531(con531),.conv532(con532),.conv533(con533),.conv534(con534),.conv535(con535),.conv536(con536),.conv537(con537),.conv538(con538),.conv539(con539),.conv540(con540),.conv541(con541),.conv542(con542),.conv543(con543),.conv544(con544),.conv545(con545),.conv546(con546),.conv547(con547),.conv548(con548),.conv549(con549),.conv550(con550),.conv551(con551),.conv552(con552),.conv553(con553),.conv554(con554),.conv555(con555),.conv556(con556),.conv557(con557),.conv558(con558),.conv559(con559),.conv560(con560),.conv561(con561),.conv562(con562),.conv563(con563),.conv564(con564),.conv565(con565),.conv566(con566),.conv567(con567),.conv568(con568),.conv569(con569),.conv570(con570),.conv571(con571),.conv572(con572),.conv573(con573),.conv574(con574),.conv575(con575),
.bias(bias),.clk(clk),.ready(readycon),.start(start));

wire [7:0] pool0;wire [7:0] pool1;wire [7:0] pool2;wire [7:0] pool3;wire [7:0] pool4;wire [7:0] pool5;wire [7:0] pool6;wire [7:0] pool7;wire [7:0] pool8;wire [7:0] pool9;wire [7:0] pool10;wire [7:0] pool11;wire [7:0] pool12;wire [7:0] pool13;wire [7:0] pool14;wire [7:0] pool15;wire [7:0] pool16;wire [7:0] pool17;wire [7:0] pool18;wire [7:0] pool19;wire [7:0] pool20;wire [7:0] pool21;wire [7:0] pool22;wire [7:0] pool23;wire [7:0] pool24;wire [7:0] pool25;wire [7:0] pool26;wire [7:0] pool27;wire [7:0] pool28;wire [7:0] pool29;wire [7:0] pool30;wire [7:0] pool31;wire [7:0] pool32;wire [7:0] pool33;wire [7:0] pool34;wire [7:0] pool35;wire [7:0] pool36;wire [7:0] pool37;wire [7:0] pool38;wire [7:0] pool39;wire [7:0] pool40;wire [7:0] pool41;wire [7:0] pool42;wire [7:0] pool43;wire [7:0] pool44;wire [7:0] pool45;wire [7:0] pool46;wire [7:0] pool47;wire [7:0] pool48;wire [7:0] pool49;wire [7:0] pool50;wire [7:0] pool51;wire [7:0] pool52;wire [7:0] pool53;wire [7:0] pool54;wire [7:0] pool55;wire [7:0] pool56;wire [7:0] pool57;wire [7:0] pool58;wire [7:0] pool59;wire [7:0] pool60;wire [7:0] pool61;wire [7:0] pool62;wire [7:0] pool63;wire [7:0] pool64;wire [7:0] pool65;wire [7:0] pool66;wire [7:0] pool67;wire [7:0] pool68;wire [7:0] pool69;wire [7:0] pool70;wire [7:0] pool71;wire [7:0] pool72;wire [7:0] pool73;wire [7:0] pool74;wire [7:0] pool75;wire [7:0] pool76;wire [7:0] pool77;wire [7:0] pool78;wire [7:0] pool79;wire [7:0] pool80;wire [7:0] pool81;wire [7:0] pool82;wire [7:0] pool83;wire [7:0] pool84;wire [7:0] pool85;wire [7:0] pool86;wire [7:0] pool87;wire [7:0] pool88;wire [7:0] pool89;wire [7:0] pool90;wire [7:0] pool91;wire [7:0] pool92;wire [7:0] pool93;wire [7:0] pool94;wire [7:0] pool95;wire [7:0] pool96;wire [7:0] pool97;wire [7:0] pool98;wire [7:0] pool99;wire [7:0] pool100;wire [7:0] pool101;wire [7:0] pool102;wire [7:0] pool103;wire [7:0] pool104;wire [7:0] pool105;wire [7:0] pool106;wire [7:0] pool107;wire [7:0] pool108;wire [7:0] pool109;wire [7:0] pool110;wire [7:0] pool111;wire [7:0] pool112;wire [7:0] pool113;wire [7:0] pool114;wire [7:0] pool115;wire [7:0] pool116;wire [7:0] pool117;wire [7:0] pool118;wire [7:0] pool119;wire [7:0] pool120;wire [7:0] pool121;wire [7:0] pool122;wire [7:0] pool123;wire [7:0] pool124;wire [7:0] pool125;wire [7:0] pool126;wire [7:0] pool127;wire [7:0] pool128;wire [7:0] pool129;wire [7:0] pool130;wire [7:0] pool131;wire [7:0] pool132;wire [7:0] pool133;wire [7:0] pool134;wire [7:0] pool135;wire [7:0] pool136;wire [7:0] pool137;wire [7:0] pool138;wire [7:0] pool139;wire [7:0] pool140;wire [7:0] pool141;wire [7:0] pool142;wire [7:0] pool143;

poolinglayer pooll1(
.in0(con0),.in1(con1),.in2(con2),.in3(con3),.in4(con4),.in5(con5),.in6(con6),.in7(con7),.in8(con8),.in9(con9),.in10(con10),.in11(con11),.in12(con12),.in13(con13),.in14(con14),.in15(con15),.in16(con16),.in17(con17),.in18(con18),.in19(con19),.in20(con20),.in21(con21),.in22(con22),.in23(con23),.in24(con24),.in25(con25),.in26(con26),.in27(con27),.in28(con28),.in29(con29),.in30(con30),.in31(con31),.in32(con32),.in33(con33),.in34(con34),.in35(con35),.in36(con36),.in37(con37),.in38(con38),.in39(con39),.in40(con40),.in41(con41),.in42(con42),.in43(con43),.in44(con44),.in45(con45),.in46(con46),.in47(con47),.in48(con48),.in49(con49),.in50(con50),.in51(con51),.in52(con52),.in53(con53),.in54(con54),.in55(con55),.in56(con56),.in57(con57),.in58(con58),.in59(con59),.in60(con60),.in61(con61),.in62(con62),.in63(con63),.in64(con64),.in65(con65),.in66(con66),.in67(con67),.in68(con68),.in69(con69),.in70(con70),.in71(con71),.in72(con72),.in73(con73),.in74(con74),.in75(con75),.in76(con76),.in77(con77),.in78(con78),.in79(con79),.in80(con80),.in81(con81),.in82(con82),.in83(con83),.in84(con84),.in85(con85),.in86(con86),.in87(con87),.in88(con88),.in89(con89),.in90(con90),.in91(con91),.in92(con92),.in93(con93),.in94(con94),.in95(con95),.in96(con96),.in97(con97),.in98(con98),.in99(con99),.in100(con100),.in101(con101),.in102(con102),.in103(con103),.in104(con104),.in105(con105),.in106(con106),.in107(con107),.in108(con108),.in109(con109),.in110(con110),.in111(con111),.in112(con112),.in113(con113),.in114(con114),.in115(con115),.in116(con116),.in117(con117),.in118(con118),.in119(con119),.in120(con120),.in121(con121),.in122(con122),.in123(con123),.in124(con124),.in125(con125),.in126(con126),.in127(con127),.in128(con128),.in129(con129),.in130(con130),.in131(con131),.in132(con132),.in133(con133),.in134(con134),.in135(con135),.in136(con136),.in137(con137),.in138(con138),.in139(con139),.in140(con140),.in141(con141),.in142(con142),.in143(con143),.in144(con144),.in145(con145),.in146(con146),.in147(con147),.in148(con148),.in149(con149),.in150(con150),.in151(con151),.in152(con152),.in153(con153),.in154(con154),.in155(con155),.in156(con156),.in157(con157),.in158(con158),.in159(con159),.in160(con160),.in161(con161),.in162(con162),.in163(con163),.in164(con164),.in165(con165),.in166(con166),.in167(con167),.in168(con168),.in169(con169),.in170(con170),.in171(con171),.in172(con172),.in173(con173),.in174(con174),.in175(con175),.in176(con176),.in177(con177),.in178(con178),.in179(con179),.in180(con180),.in181(con181),.in182(con182),.in183(con183),.in184(con184),.in185(con185),.in186(con186),.in187(con187),.in188(con188),.in189(con189),.in190(con190),.in191(con191),.in192(con192),.in193(con193),.in194(con194),.in195(con195),.in196(con196),.in197(con197),.in198(con198),.in199(con199),.in200(con200),.in201(con201),.in202(con202),.in203(con203),.in204(con204),.in205(con205),.in206(con206),.in207(con207),.in208(con208),.in209(con209),.in210(con210),.in211(con211),.in212(con212),.in213(con213),.in214(con214),.in215(con215),.in216(con216),.in217(con217),.in218(con218),.in219(con219),.in220(con220),.in221(con221),.in222(con222),.in223(con223),.in224(con224),.in225(con225),.in226(con226),.in227(con227),.in228(con228),.in229(con229),.in230(con230),.in231(con231),.in232(con232),.in233(con233),.in234(con234),.in235(con235),.in236(con236),.in237(con237),.in238(con238),.in239(con239),.in240(con240),.in241(con241),.in242(con242),.in243(con243),.in244(con244),.in245(con245),.in246(con246),.in247(con247),.in248(con248),.in249(con249),.in250(con250),.in251(con251),.in252(con252),.in253(con253),.in254(con254),.in255(con255),.in256(con256),.in257(con257),.in258(con258),.in259(con259),.in260(con260),.in261(con261),.in262(con262),.in263(con263),.in264(con264),.in265(con265),.in266(con266),.in267(con267),.in268(con268),.in269(con269),.in270(con270),.in271(con271),.in272(con272),.in273(con273),.in274(con274),.in275(con275),.in276(con276),.in277(con277),.in278(con278),.in279(con279),.in280(con280),.in281(con281),.in282(con282),.in283(con283),.in284(con284),.in285(con285),.in286(con286),.in287(con287),.in288(con288),.in289(con289),.in290(con290),.in291(con291),.in292(con292),.in293(con293),.in294(con294),.in295(con295),.in296(con296),.in297(con297),.in298(con298),.in299(con299),.in300(con300),.in301(con301),.in302(con302),.in303(con303),.in304(con304),.in305(con305),.in306(con306),.in307(con307),.in308(con308),.in309(con309),.in310(con310),.in311(con311),.in312(con312),.in313(con313),.in314(con314),.in315(con315),.in316(con316),.in317(con317),.in318(con318),.in319(con319),.in320(con320),.in321(con321),.in322(con322),.in323(con323),.in324(con324),.in325(con325),.in326(con326),.in327(con327),.in328(con328),.in329(con329),.in330(con330),.in331(con331),.in332(con332),.in333(con333),.in334(con334),.in335(con335),.in336(con336),.in337(con337),.in338(con338),.in339(con339),.in340(con340),.in341(con341),.in342(con342),.in343(con343),.in344(con344),.in345(con345),.in346(con346),.in347(con347),.in348(con348),.in349(con349),.in350(con350),.in351(con351),.in352(con352),.in353(con353),.in354(con354),.in355(con355),.in356(con356),.in357(con357),.in358(con358),.in359(con359),.in360(con360),.in361(con361),.in362(con362),.in363(con363),.in364(con364),.in365(con365),.in366(con366),.in367(con367),.in368(con368),.in369(con369),.in370(con370),.in371(con371),.in372(con372),.in373(con373),.in374(con374),.in375(con375),.in376(con376),.in377(con377),.in378(con378),.in379(con379),.in380(con380),.in381(con381),.in382(con382),.in383(con383),.in384(con384),.in385(con385),.in386(con386),.in387(con387),.in388(con388),.in389(con389),.in390(con390),.in391(con391),.in392(con392),.in393(con393),.in394(con394),.in395(con395),.in396(con396),.in397(con397),.in398(con398),.in399(con399),.in400(con400),.in401(con401),.in402(con402),.in403(con403),.in404(con404),.in405(con405),.in406(con406),.in407(con407),.in408(con408),.in409(con409),.in410(con410),.in411(con411),.in412(con412),.in413(con413),.in414(con414),.in415(con415),.in416(con416),.in417(con417),.in418(con418),.in419(con419),.in420(con420),.in421(con421),.in422(con422),.in423(con423),.in424(con424),.in425(con425),.in426(con426),.in427(con427),.in428(con428),.in429(con429),.in430(con430),.in431(con431),.in432(con432),.in433(con433),.in434(con434),.in435(con435),.in436(con436),.in437(con437),.in438(con438),.in439(con439),.in440(con440),.in441(con441),.in442(con442),.in443(con443),.in444(con444),.in445(con445),.in446(con446),.in447(con447),.in448(con448),.in449(con449),.in450(con450),.in451(con451),.in452(con452),.in453(con453),.in454(con454),.in455(con455),.in456(con456),.in457(con457),.in458(con458),.in459(con459),.in460(con460),.in461(con461),.in462(con462),.in463(con463),.in464(con464),.in465(con465),.in466(con466),.in467(con467),.in468(con468),.in469(con469),.in470(con470),.in471(con471),.in472(con472),.in473(con473),.in474(con474),.in475(con475),.in476(con476),.in477(con477),.in478(con478),.in479(con479),.in480(con480),.in481(con481),.in482(con482),.in483(con483),.in484(con484),.in485(con485),.in486(con486),.in487(con487),.in488(con488),.in489(con489),.in490(con490),.in491(con491),.in492(con492),.in493(con493),.in494(con494),.in495(con495),.in496(con496),.in497(con497),.in498(con498),.in499(con499),.in500(con500),.in501(con501),.in502(con502),.in503(con503),.in504(con504),.in505(con505),.in506(con506),.in507(con507),.in508(con508),.in509(con509),.in510(con510),.in511(con511),.in512(con512),.in513(con513),.in514(con514),.in515(con515),.in516(con516),.in517(con517),.in518(con518),.in519(con519),.in520(con520),.in521(con521),.in522(con522),.in523(con523),.in524(con524),.in525(con525),.in526(con526),.in527(con527),.in528(con528),.in529(con529),.in530(con530),.in531(con531),.in532(con532),.in533(con533),.in534(con534),.in535(con535),.in536(con536),.in537(con537),.in538(con538),.in539(con539),.in540(con540),.in541(con541),.in542(con542),.in543(con543),.in544(con544),.in545(con545),.in546(con546),.in547(con547),.in548(con548),.in549(con549),.in550(con550),.in551(con551),.in552(con552),.in553(con553),.in554(con554),.in555(con555),.in556(con556),.in557(con557),.in558(con558),.in559(con559),.in560(con560),.in561(con561),.in562(con562),.in563(con563),.in564(con564),.in565(con565),.in566(con566),.in567(con567),.in568(con568),.in569(con569),.in570(con570),.in571(con571),.in572(con572),.in573(con573),.in574(con574),.in575(con575),
.out0(pool0),.out1(pool1),.out2(pool2),.out3(pool3),.out4(pool4),.out5(pool5),.out6(pool6),.out7(pool7),.out8(pool8),.out9(pool9),.out10(pool10),.out11(pool11),.out12(pool12),.out13(pool13),.out14(pool14),.out15(pool15),.out16(pool16),.out17(pool17),.out18(pool18),.out19(pool19),.out20(pool20),.out21(pool21),.out22(pool22),.out23(pool23),.out24(pool24),.out25(pool25),.out26(pool26),.out27(pool27),.out28(pool28),.out29(pool29),.out30(pool30),.out31(pool31),.out32(pool32),.out33(pool33),.out34(pool34),.out35(pool35),.out36(pool36),.out37(pool37),.out38(pool38),.out39(pool39),.out40(pool40),.out41(pool41),.out42(pool42),.out43(pool43),.out44(pool44),.out45(pool45),.out46(pool46),.out47(pool47),.out48(pool48),.out49(pool49),.out50(pool50),.out51(pool51),.out52(pool52),.out53(pool53),.out54(pool54),.out55(pool55),.out56(pool56),.out57(pool57),.out58(pool58),.out59(pool59),.out60(pool60),.out61(pool61),.out62(pool62),.out63(pool63),.out64(pool64),.out65(pool65),.out66(pool66),.out67(pool67),.out68(pool68),.out69(pool69),.out70(pool70),.out71(pool71),.out72(pool72),.out73(pool73),.out74(pool74),.out75(pool75),.out76(pool76),.out77(pool77),.out78(pool78),.out79(pool79),.out80(pool80),.out81(pool81),.out82(pool82),.out83(pool83),.out84(pool84),.out85(pool85),.out86(pool86),.out87(pool87),.out88(pool88),.out89(pool89),.out90(pool90),.out91(pool91),.out92(pool92),.out93(pool93),.out94(pool94),.out95(pool95),.out96(pool96),.out97(pool97),.out98(pool98),.out99(pool99),.out100(pool100),.out101(pool101),.out102(pool102),.out103(pool103),.out104(pool104),.out105(pool105),.out106(pool106),.out107(pool107),.out108(pool108),.out109(pool109),.out110(pool110),.out111(pool111),.out112(pool112),.out113(pool113),.out114(pool114),.out115(pool115),.out116(pool116),.out117(pool117),.out118(pool118),.out119(pool119),.out120(pool120),.out121(pool121),.out122(pool122),.out123(pool123),.out124(pool124),.out125(pool125),.out126(pool126),.out127(pool127),.out128(pool128),.out129(pool129),.out130(pool130),.out131(pool131),.out132(pool132),.out133(pool133),.out134(pool134),.out135(pool135),.out136(pool136),.out137(pool137),.out138(pool138),.out139(pool139),.out140(pool140),.out141(pool141),.out142(pool142),.out143(pool143),
.clk(clk),.ready(readypool),.start(readycon));



FullyConnected F1(.weight0(weight2l0),.weight1(weight2l1),.weight2(weight2l2),.weight3(weight2l3),.weight4(weight2l4),.weight5(weight2l5),.weight6(weight2l6),.weight7(weight2l7),.weight8(weight2l8),.weight9(weight2l9),.weight10(weight2l10),.weight11(weight2l11),.weight12(weight2l12),.weight13(weight2l13),.weight14(weight2l14),.weight15(weight2l15),.weight16(weight2l16),.weight17(weight2l17),.weight18(weight2l18),.weight19(weight2l19),.weight20(weight2l20),.weight21(weight2l21),.weight22(weight2l22),.weight23(weight2l23),.weight24(weight2l24),.weight25(weight2l25),.weight26(weight2l26),.weight27(weight2l27),.weight28(weight2l28),.weight29(weight2l29),.weight30(weight2l30),.weight31(weight2l31),.weight32(weight2l32),.weight33(weight2l33),.weight34(weight2l34),.weight35(weight2l35),.weight36(weight2l36),.weight37(weight2l37),.weight38(weight2l38),.weight39(weight2l39),.weight40(weight2l40),.weight41(weight2l41),.weight42(weight2l42),.weight43(weight2l43),.weight44(weight2l44),.weight45(weight2l45),.weight46(weight2l46),.weight47(weight2l47),.weight48(weight2l48),.weight49(weight2l49),.weight50(weight2l50),.weight51(weight2l51),.weight52(weight2l52),.weight53(weight2l53),.weight54(weight2l54),.weight55(weight2l55),.weight56(weight2l56),.weight57(weight2l57),.weight58(weight2l58),.weight59(weight2l59),.weight60(weight2l60),.weight61(weight2l61),.weight62(weight2l62),.weight63(weight2l63),.weight64(weight2l64),.weight65(weight2l65),.weight66(weight2l66),.weight67(weight2l67),.weight68(weight2l68),.weight69(weight2l69),.weight70(weight2l70),.weight71(weight2l71),.weight72(weight2l72),.weight73(weight2l73),.weight74(weight2l74),.weight75(weight2l75),.weight76(weight2l76),.weight77(weight2l77),.weight78(weight2l78),.weight79(weight2l79),.weight80(weight2l80),.weight81(weight2l81),.weight82(weight2l82),.weight83(weight2l83),.weight84(weight2l84),.weight85(weight2l85),.weight86(weight2l86),.weight87(weight2l87),.weight88(weight2l88),.weight89(weight2l89),.weight90(weight2l90),.weight91(weight2l91),.weight92(weight2l92),.weight93(weight2l93),.weight94(weight2l94),.weight95(weight2l95),.weight96(weight2l96),.weight97(weight2l97),.weight98(weight2l98),.weight99(weight2l99),.weight100(weight2l100),.weight101(weight2l101),.weight102(weight2l102),.weight103(weight2l103),.weight104(weight2l104),.weight105(weight2l105),.weight106(weight2l106),.weight107(weight2l107),.weight108(weight2l108),.weight109(weight2l109),.weight110(weight2l110),.weight111(weight2l111),.weight112(weight2l112),.weight113(weight2l113),.weight114(weight2l114),.weight115(weight2l115),.weight116(weight2l116),.weight117(weight2l117),.weight118(weight2l118),.weight119(weight2l119),.weight120(weight2l120),.weight121(weight2l121),.weight122(weight2l122),.weight123(weight2l123),.weight124(weight2l124),.weight125(weight2l125),.weight126(weight2l126),.weight127(weight2l127),.weight128(weight2l128),.weight129(weight2l129),.weight130(weight2l130),.weight131(weight2l131),.weight132(weight2l132),.weight133(weight2l133),.weight134(weight2l134),.weight135(weight2l135),.weight136(weight2l136),.weight137(weight2l137),.weight138(weight2l138),.weight139(weight2l139),.weight140(weight2l140),.weight141(weight2l141),.weight142(weight2l142),.weight143(weight2l143),
.in0(pool0),.in1(pool1),.in2(pool2),.in3(pool3),.in4(pool4),.in5(pool5),.in6(pool6),.in7(pool7),.in8(pool8),.in9(pool9),.in10(pool10),.in11(pool11),.in12(pool12),.in13(pool13),.in14(pool14),.in15(pool15),.in16(pool16),.in17(pool17),.in18(pool18),.in19(pool19),.in20(pool20),.in21(pool21),.in22(pool22),.in23(pool23),.in24(pool24),.in25(pool25),.in26(pool26),.in27(pool27),.in28(pool28),.in29(pool29),.in30(pool30),.in31(pool31),.in32(pool32),.in33(pool33),.in34(pool34),.in35(pool35),.in36(pool36),.in37(pool37),.in38(pool38),.in39(pool39),.in40(pool40),.in41(pool41),.in42(pool42),.in43(pool43),.in44(pool44),.in45(pool45),.in46(pool46),.in47(pool47),.in48(pool48),.in49(pool49),.in50(pool50),.in51(pool51),.in52(pool52),.in53(pool53),.in54(pool54),.in55(pool55),.in56(pool56),.in57(pool57),.in58(pool58),.in59(pool59),.in60(pool60),.in61(pool61),.in62(pool62),.in63(pool63),.in64(pool64),.in65(pool65),.in66(pool66),.in67(pool67),.in68(pool68),.in69(pool69),.in70(pool70),.in71(pool71),.in72(pool72),.in73(pool73),.in74(pool74),.in75(pool75),.in76(pool76),.in77(pool77),.in78(pool78),.in79(pool79),.in80(pool80),.in81(pool81),.in82(pool82),.in83(pool83),.in84(pool84),.in85(pool85),.in86(pool86),.in87(pool87),.in88(pool88),.in89(pool89),.in90(pool90),.in91(pool91),.in92(pool92),.in93(pool93),.in94(pool94),.in95(pool95),.in96(pool96),.in97(pool97),.in98(pool98),.in99(pool99),.in100(pool100),.in101(pool101),.in102(pool102),.in103(pool103),.in104(pool104),.in105(pool105),.in106(pool106),.in107(pool107),.in108(pool108),.in109(pool109),.in110(pool110),.in111(pool111),.in112(pool112),.in113(pool113),.in114(pool114),.in115(pool115),.in116(pool116),.in117(pool117),.in118(pool118),.in119(pool119),.in120(pool120),.in121(pool121),.in122(pool122),.in123(pool123),.in124(pool124),.in125(pool125),.in126(pool126),.in127(pool127),.in128(pool128),.in129(pool129),.in130(pool130),.in131(pool131),.in132(pool132),.in133(pool133),.in134(pool134),.in135(pool135),.in136(pool136),.in137(pool137),.in138(pool138),.in139(pool139),.in140(pool140),.in141(pool141),.in142(pool142),.in143(pool143),
.clk(clk),.start(readypool),.ready(ready),.out(out));

endmodule
