`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    09:53:34 11/07/2017 
// Design Name: 
// Module Name:    FullyConnected 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module FullyConnected(
weight0,weight1,weight2,weight3,weight4,weight5,weight6,weight7,weight8,weight9,weight10,weight11,weight12,weight13,weight14,weight15,weight16,weight17,weight18,weight19,weight20,weight21,weight22,weight23,weight24,weight25,weight26,weight27,weight28,weight29,weight30,weight31,weight32,weight33,weight34,weight35,weight36,weight37,weight38,weight39,weight40,weight41,weight42,weight43,weight44,weight45,weight46,weight47,weight48,weight49,weight50,weight51,weight52,weight53,weight54,weight55,weight56,weight57,weight58,weight59,weight60,weight61,weight62,weight63,weight64,weight65,weight66,weight67,weight68,weight69,weight70,weight71,weight72,weight73,weight74,weight75,weight76,weight77,weight78,weight79,weight80,weight81,weight82,weight83,weight84,weight85,weight86,weight87,weight88,weight89,weight90,weight91,weight92,weight93,weight94,weight95,weight96,weight97,weight98,weight99,weight100,weight101,weight102,weight103,weight104,weight105,weight106,weight107,weight108,weight109,weight110,weight111,weight112,weight113,weight114,weight115,weight116,weight117,weight118,weight119,weight120,weight121,weight122,weight123,weight124,weight125,weight126,weight127,weight128,weight129,weight130,weight131,weight132,weight133,weight134,weight135,weight136,weight137,weight138,weight139,weight140,weight141,weight142,weight143,
in0,in1,in2,in3,in4,in5,in6,in7,in8,in9,in10,in11,in12,in13,in14,in15,in16,in17,in18,in19,in20,in21,in22,in23,in24,in25,in26,in27,in28,in29,in30,in31,in32,in33,in34,in35,in36,in37,in38,in39,in40,in41,in42,in43,in44,in45,in46,in47,in48,in49,in50,in51,in52,in53,in54,in55,in56,in57,in58,in59,in60,in61,in62,in63,in64,in65,in66,in67,in68,in69,in70,in71,in72,in73,in74,in75,in76,in77,in78,in79,in80,in81,in82,in83,in84,in85,in86,in87,in88,in89,in90,in91,in92,in93,in94,in95,in96,in97,in98,in99,in100,in101,in102,in103,in104,in105,in106,in107,in108,in109,in110,in111,in112,in113,in114,in115,in116,in117,in118,in119,in120,in121,in122,in123,in124,in125,in126,in127,in128,in129,in130,in131,in132,in133,in134,in135,in136,in137,in138,in139,in140,in141,in142,in143,
clk,start,out,ready);

input start;
input clk;
output ready;
reg ready;
output [7:0] out;
input [7:0] in0;
input [7:0] in1;
input [7:0] in2;
input [7:0] in3;
input [7:0] in4;
input [7:0] in5;
input [7:0] in6;
input [7:0] in7;
input [7:0] in8;
input [7:0] in9;
input [7:0] in10;
input [7:0] in11;
input [7:0] in12;
input [7:0] in13;
input [7:0] in14;
input [7:0] in15;
input [7:0] in16;
input [7:0] in17;
input [7:0] in18;
input [7:0] in19;
input [7:0] in20;
input [7:0] in21;
input [7:0] in22;
input [7:0] in23;
input [7:0] in24;
input [7:0] in25;
input [7:0] in26;
input [7:0] in27;
input [7:0] in28;
input [7:0] in29;
input [7:0] in30;
input [7:0] in31;
input [7:0] in32;
input [7:0] in33;
input [7:0] in34;
input [7:0] in35;
input [7:0] in36;
input [7:0] in37;
input [7:0] in38;
input [7:0] in39;
input [7:0] in40;
input [7:0] in41;
input [7:0] in42;
input [7:0] in43;
input [7:0] in44;
input [7:0] in45;
input [7:0] in46;
input [7:0] in47;
input [7:0] in48;
input [7:0] in49;
input [7:0] in50;
input [7:0] in51;
input [7:0] in52;
input [7:0] in53;
input [7:0] in54;
input [7:0] in55;
input [7:0] in56;
input [7:0] in57;
input [7:0] in58;
input [7:0] in59;
input [7:0] in60;
input [7:0] in61;
input [7:0] in62;
input [7:0] in63;
input [7:0] in64;
input [7:0] in65;
input [7:0] in66;
input [7:0] in67;
input [7:0] in68;
input [7:0] in69;
input [7:0] in70;
input [7:0] in71;
input [7:0] in72;
input [7:0] in73;
input [7:0] in74;
input [7:0] in75;
input [7:0] in76;
input [7:0] in77;
input [7:0] in78;
input [7:0] in79;
input [7:0] in80;
input [7:0] in81;
input [7:0] in82;
input [7:0] in83;
input [7:0] in84;
input [7:0] in85;
input [7:0] in86;
input [7:0] in87;
input [7:0] in88;
input [7:0] in89;
input [7:0] in90;
input [7:0] in91;
input [7:0] in92;
input [7:0] in93;
input [7:0] in94;
input [7:0] in95;
input [7:0] in96;
input [7:0] in97;
input [7:0] in98;
input [7:0] in99;
input [7:0] in100;
input [7:0] in101;
input [7:0] in102;
input [7:0] in103;
input [7:0] in104;
input [7:0] in105;
input [7:0] in106;
input [7:0] in107;
input [7:0] in108;
input [7:0] in109;
input [7:0] in110;
input [7:0] in111;
input [7:0] in112;
input [7:0] in113;
input [7:0] in114;
input [7:0] in115;
input [7:0] in116;
input [7:0] in117;
input [7:0] in118;
input [7:0] in119;
input [7:0] in120;
input [7:0] in121;
input [7:0] in122;
input [7:0] in123;
input [7:0] in124;
input [7:0] in125;
input [7:0] in126;
input [7:0] in127;
input [7:0] in128;
input [7:0] in129;
input [7:0] in130;
input [7:0] in131;
input [7:0] in132;
input [7:0] in133;
input [7:0] in134;
input [7:0] in135;
input [7:0] in136;
input [7:0] in137;
input [7:0] in138;
input [7:0] in139;
input [7:0] in140;
input [7:0] in141;
input [7:0] in142;
input [7:0] in143;

 input [7:0] weight0;
input [7:0] weight1;
input [7:0] weight2;
input [7:0] weight3;
input [7:0] weight4;
input [7:0] weight5;
input [7:0] weight6;
input [7:0] weight7;
input [7:0] weight8;
input [7:0] weight9;
input [7:0] weight10;
input [7:0] weight11;
input [7:0] weight12;
input [7:0] weight13;
input [7:0] weight14;
input [7:0] weight15;
input [7:0] weight16;
input [7:0] weight17;
input [7:0] weight18;
input [7:0] weight19;
input [7:0] weight20;
input [7:0] weight21;
input [7:0] weight22;
input [7:0] weight23;
input [7:0] weight24;
input [7:0] weight25;
input [7:0] weight26;
input [7:0] weight27;
input [7:0] weight28;
input [7:0] weight29;
input [7:0] weight30;
input [7:0] weight31;
input [7:0] weight32;
input [7:0] weight33;
input [7:0] weight34;
input [7:0] weight35;
input [7:0] weight36;
input [7:0] weight37;
input [7:0] weight38;
input [7:0] weight39;
input [7:0] weight40;
input [7:0] weight41;
input [7:0] weight42;
input [7:0] weight43;
input [7:0] weight44;
input [7:0] weight45;
input [7:0] weight46;
input [7:0] weight47;
input [7:0] weight48;
input [7:0] weight49;
input [7:0] weight50;
input [7:0] weight51;
input [7:0] weight52;
input [7:0] weight53;
input [7:0] weight54;
input [7:0] weight55;
input [7:0] weight56;
input [7:0] weight57;
input [7:0] weight58;
input [7:0] weight59;
input [7:0] weight60;
input [7:0] weight61;
input [7:0] weight62;
input [7:0] weight63;
input [7:0] weight64;
input [7:0] weight65;
input [7:0] weight66;
input [7:0] weight67;
input [7:0] weight68;
input [7:0] weight69;
input [7:0] weight70;
input [7:0] weight71;
input [7:0] weight72;
input [7:0] weight73;
input [7:0] weight74;
input [7:0] weight75;
input [7:0] weight76;
input [7:0] weight77;
input [7:0] weight78;
input [7:0] weight79;
input [7:0] weight80;
input [7:0] weight81;
input [7:0] weight82;
input [7:0] weight83;
input [7:0] weight84;
input [7:0] weight85;
input [7:0] weight86;
input [7:0] weight87;
input [7:0] weight88;
input [7:0] weight89;
input [7:0] weight90;
input [7:0] weight91;
input [7:0] weight92;
input [7:0] weight93;
input [7:0] weight94;
input [7:0] weight95;
input [7:0] weight96;
input [7:0] weight97;
input [7:0] weight98;
input [7:0] weight99;
input [7:0] weight100;
input [7:0] weight101;
input [7:0] weight102;
input [7:0] weight103;
input [7:0] weight104;
input [7:0] weight105;
input [7:0] weight106;
input [7:0] weight107;
input [7:0] weight108;
input [7:0] weight109;
input [7:0] weight110;
input [7:0] weight111;
input [7:0] weight112;
input [7:0] weight113;
input [7:0] weight114;
input [7:0] weight115;
input [7:0] weight116;
input [7:0] weight117;
input [7:0] weight118;
input [7:0] weight119;
input [7:0] weight120;
input [7:0] weight121;
input [7:0] weight122;
input [7:0] weight123;
input [7:0] weight124;
input [7:0] weight125;
input [7:0] weight126;
input [7:0] weight127;
input [7:0] weight128;
input [7:0] weight129;
input [7:0] weight130;
input [7:0] weight131;
input [7:0] weight132;
input [7:0] weight133;
input [7:0] weight134;
input [7:0] weight135;
input [7:0] weight136;
input [7:0] weight137;
input [7:0] weight138;
input [7:0] weight139;
input [7:0] weight140;
input [7:0] weight141;
input [7:0] weight142;
input [7:0] weight143;



wire [7:0] mux0;
wire [7:0] mux1;
wire [7:0] mux2;
wire [7:0] mux3;
wire [7:0] mux4;
wire [7:0] mux5;
wire [7:0] mux6;
wire [7:0] mux7;
wire [7:0] mux8;
wire [7:0] mux9;
wire [7:0] mux10;
wire [7:0] mux11;
wire [7:0] mux12;
wire [7:0] mux13;
wire [7:0] mux14;
wire [7:0] mux15;
wire [7:0] mux16;
wire [7:0] mux17;
wire [7:0] mux18;
wire [7:0] mux19;
wire [7:0] mux20;
wire [7:0] mux21;
wire [7:0] mux22;
wire [7:0] mux23;
wire [7:0] mux24;
wire [7:0] mux25;
wire [7:0] mux26;
wire [7:0] mux27;
wire [7:0] mux28;
wire [7:0] mux29;
wire [7:0] mux30;
wire [7:0] mux31;
wire [7:0] mux32;
wire [7:0] mux33;
wire [7:0] mux34;
wire [7:0] mux35;

 wire [7:0] mulo0;
wire [7:0] mulo1;
wire [7:0] mulo2;
wire [7:0] mulo3;
wire [7:0] mulo4;
wire [7:0] mulo5;
wire [7:0] mulo6;
wire [7:0] mulo7;
wire [7:0] mulo8;
wire [7:0] mulo9;
wire [7:0] mulo10;
wire [7:0] mulo11;
wire [7:0] mulo12;
wire [7:0] mulo13;
wire [7:0] mulo14;
wire [7:0] mulo15;
wire [7:0] mulo16;
wire [7:0] mulo17;
wire [7:0] mulo18;
wire [7:0] mulo19;
wire [7:0] mulo20;
wire [7:0] mulo21;
wire [7:0] mulo22;
wire [7:0] mulo23;
wire [7:0] mulo24;
wire [7:0] mulo25;
wire [7:0] mulo26;
wire [7:0] mulo27;
wire [7:0] mulo28;
wire [7:0] mulo29;
wire [7:0] mulo30;
wire [7:0] mulo31;
wire [7:0] mulo32;
wire [7:0] mulo33;
wire [7:0] mulo34;
wire [7:0] mulo35;

 wire [7:0] muxo0;
wire [7:0] muxo1;
wire [7:0] muxo2;
wire [7:0] muxo3;
wire [7:0] muxo4;
wire [7:0] muxo5;
wire [7:0] muxo6;
wire [7:0] muxo7;
wire [7:0] muxo8;
wire [7:0] muxo9;
wire [7:0] muxo10;
wire [7:0] muxo11;
wire [7:0] muxo12;
wire [7:0] muxo13;
wire [7:0] muxo14;
wire [7:0] muxo15;
wire [7:0] muxo16;
wire [7:0] muxo17;
wire [7:0] muxo18;
wire [7:0] muxo19;
wire [7:0] muxo20;
wire [7:0] muxo21;
wire [7:0] muxo22;
wire [7:0] muxo23;
wire [7:0] muxo24;
wire [7:0] muxo25;
wire [7:0] muxo26;
wire [7:0] muxo27;
wire [7:0] muxo28;
wire [7:0] muxo29;
wire [7:0] muxo30;
wire [7:0] muxo31;
wire [7:0] muxo32;
wire [7:0] muxo33;
wire [7:0] muxo34;
wire [7:0] muxo35;
wire [7:0] muxo36;
wire [7:0] muxo37;
wire [7:0] muxo38;
wire [7:0] muxo39;
wire [7:0] muxo40;
wire [7:0] muxo41;
wire [7:0] muxo42;
wire [7:0] muxo43;
wire [7:0] muxo44;
wire [7:0] muxo45;
wire [7:0] muxo46;
wire [7:0] muxo47;
wire [7:0] muxo48;
wire [7:0] muxo49;
wire [7:0] muxo50;
wire [7:0] muxo51;
wire [7:0] muxo52;
wire [7:0] muxo53;
wire [7:0] muxo54;
wire [7:0] muxo55;
wire [7:0] muxo56;
wire [7:0] muxo57;
wire [7:0] muxo58;
wire [7:0] muxo59;
wire [7:0] muxo60;
wire [7:0] muxo61;
wire [7:0] muxo62;
wire [7:0] muxo63;
wire [7:0] muxo64;
wire [7:0] muxo65;
wire [7:0] muxo66;
wire [7:0] muxo67;
wire [7:0] muxo68;
wire [7:0] muxo69;
wire [7:0] muxo70;
wire [7:0] muxo71;
wire [7:0] muxo72;
wire [7:0] muxo73;
wire [7:0] muxo74;
wire [7:0] muxo75;
wire [7:0] muxo76;
wire [7:0] muxo77;
wire [7:0] muxo78;
wire [7:0] muxo79;
wire [7:0] muxo80;
wire [7:0] muxo81;
wire [7:0] muxo82;
wire [7:0] muxo83;
wire [7:0] muxo84;
wire [7:0] muxo85;
wire [7:0] muxo86;
wire [7:0] muxo87;
wire [7:0] muxo88;
wire [7:0] muxo89;
wire [7:0] muxo90;
wire [7:0] muxo91;
wire [7:0] muxo92;
wire [7:0] muxo93;
wire [7:0] muxo94;
wire [7:0] muxo95;
wire [7:0] muxo96;
wire [7:0] muxo97;
wire [7:0] muxo98;
wire [7:0] muxo99;
wire [7:0] muxo100;
wire [7:0] muxo101;
wire [7:0] muxo102;
wire [7:0] muxo103;
wire [7:0] muxo104;
wire [7:0] muxo105;
wire [7:0] muxo106;
wire [7:0] muxo107;
wire [7:0] muxo108;
wire [7:0] muxo109;
wire [7:0] muxo110;
wire [7:0] muxo111;
wire [7:0] muxo112;
wire [7:0] muxo113;
wire [7:0] muxo114;
wire [7:0] muxo115;
wire [7:0] muxo116;
wire [7:0] muxo117;
wire [7:0] muxo118;
wire [7:0] muxo119;
wire [7:0] muxo120;
wire [7:0] muxo121;
wire [7:0] muxo122;
wire [7:0] muxo123;
wire [7:0] muxo124;
wire [7:0] muxo125;
wire [7:0] muxo126;
wire [7:0] muxo127;
wire [7:0] muxo128;
wire [7:0] muxo129;
wire [7:0] muxo130;
wire [7:0] muxo131;
wire [7:0] muxo132;
wire [7:0] muxo133;
wire [7:0] muxo134;
wire [7:0] muxo135;
wire [7:0] muxo136;
wire [7:0] muxo137;
wire [7:0] muxo138;
wire [7:0] muxo139;
wire [7:0] muxo140;
wire [7:0] muxo141;
wire [7:0] muxo142;
wire [7:0] muxo143;


 wire [7:0] muxw0;
wire [7:0] muxw1;
wire [7:0] muxw2;
wire [7:0] muxw3;
wire [7:0] muxw4;
wire [7:0] muxw5;
wire [7:0] muxw6;
wire [7:0] muxw7;
wire [7:0] muxw8;
wire [7:0] muxw9;
wire [7:0] muxw10;
wire [7:0] muxw11;
wire [7:0] muxw12;
wire [7:0] muxw13;
wire [7:0] muxw14;
wire [7:0] muxw15;
wire [7:0] muxw16;
wire [7:0] muxw17;
wire [7:0] muxw18;
wire [7:0] muxw19;
wire [7:0] muxw20;
wire [7:0] muxw21;
wire [7:0] muxw22;
wire [7:0] muxw23;
wire [7:0] muxw24;
wire [7:0] muxw25;
wire [7:0] muxw26;
wire [7:0] muxw27;
wire [7:0] muxw28;
wire [7:0] muxw29;
wire [7:0] muxw30;
wire [7:0] muxw31;
wire [7:0] muxw32;
wire [7:0] muxw33;
wire [7:0] muxw34;
wire [7:0] muxw35;


reg [3:0] cs;

assign out = outreg;


mux42 mux42fi0(.a(in0),.b(in36),.c(in72),.d(in108),.sel(cs[1:0]),.out(mux0));
mux42 mux42fi1(.a(in1),.b(in37),.c(in73),.d(in109),.sel(cs[1:0]),.out(mux1));
mux42 mux42fi2(.a(in2),.b(in38),.c(in74),.d(in110),.sel(cs[1:0]),.out(mux2));
mux42 mux42fi3(.a(in3),.b(in39),.c(in75),.d(in111),.sel(cs[1:0]),.out(mux3));
mux42 mux42fi4(.a(in4),.b(in40),.c(in76),.d(in112),.sel(cs[1:0]),.out(mux4));
mux42 mux42fi5(.a(in5),.b(in41),.c(in77),.d(in113),.sel(cs[1:0]),.out(mux5));
mux42 mux42fi6(.a(in6),.b(in42),.c(in78),.d(in114),.sel(cs[1:0]),.out(mux6));
mux42 mux42fi7(.a(in7),.b(in43),.c(in79),.d(in115),.sel(cs[1:0]),.out(mux7));
mux42 mux42fi8(.a(in8),.b(in44),.c(in80),.d(in116),.sel(cs[1:0]),.out(mux8));
mux42 mux42fi9(.a(in9),.b(in45),.c(in81),.d(in117),.sel(cs[1:0]),.out(mux9));
mux42 mux42fi10(.a(in10),.b(in46),.c(in82),.d(in118),.sel(cs[1:0]),.out(mux10));
mux42 mux42fi11(.a(in11),.b(in47),.c(in83),.d(in119),.sel(cs[1:0]),.out(mux11));
mux42 mux42fi12(.a(in12),.b(in48),.c(in84),.d(in120),.sel(cs[1:0]),.out(mux12));
mux42 mux42fi13(.a(in13),.b(in49),.c(in85),.d(in121),.sel(cs[1:0]),.out(mux13));
mux42 mux42fi14(.a(in14),.b(in50),.c(in86),.d(in122),.sel(cs[1:0]),.out(mux14));
mux42 mux42fi15(.a(in15),.b(in51),.c(in87),.d(in123),.sel(cs[1:0]),.out(mux15));
mux42 mux42fi16(.a(in16),.b(in52),.c(in88),.d(in124),.sel(cs[1:0]),.out(mux16));
mux42 mux42fi17(.a(in17),.b(in53),.c(in89),.d(in125),.sel(cs[1:0]),.out(mux17));
mux42 mux42fi18(.a(in18),.b(in54),.c(in90),.d(in126),.sel(cs[1:0]),.out(mux18));
mux42 mux42fi19(.a(in19),.b(in55),.c(in91),.d(in127),.sel(cs[1:0]),.out(mux19));
mux42 mux42fi20(.a(in20),.b(in56),.c(in92),.d(in128),.sel(cs[1:0]),.out(mux20));
mux42 mux42fi21(.a(in21),.b(in57),.c(in93),.d(in129),.sel(cs[1:0]),.out(mux21));
mux42 mux42fi22(.a(in22),.b(in58),.c(in94),.d(in130),.sel(cs[1:0]),.out(mux22));
mux42 mux42fi23(.a(in23),.b(in59),.c(in95),.d(in131),.sel(cs[1:0]),.out(mux23));
mux42 mux42fi24(.a(in24),.b(in60),.c(in96),.d(in132),.sel(cs[1:0]),.out(mux24));
mux42 mux42fi25(.a(in25),.b(in61),.c(in97),.d(in133),.sel(cs[1:0]),.out(mux25));
mux42 mux42fi26(.a(in26),.b(in62),.c(in98),.d(in134),.sel(cs[1:0]),.out(mux26));
mux42 mux42fi27(.a(in27),.b(in63),.c(in99),.d(in135),.sel(cs[1:0]),.out(mux27));
mux42 mux42fi28(.a(in28),.b(in64),.c(in100),.d(in136),.sel(cs[1:0]),.out(mux28));
mux42 mux42fi29(.a(in29),.b(in65),.c(in101),.d(in137),.sel(cs[1:0]),.out(mux29));
mux42 mux42fi30(.a(in30),.b(in66),.c(in102),.d(in138),.sel(cs[1:0]),.out(mux30));
mux42 mux42fi31(.a(in31),.b(in67),.c(in103),.d(in139),.sel(cs[1:0]),.out(mux31));
mux42 mux42fi32(.a(in32),.b(in68),.c(in104),.d(in140),.sel(cs[1:0]),.out(mux32));
mux42 mux42fi33(.a(in33),.b(in69),.c(in105),.d(in141),.sel(cs[1:0]),.out(mux33));
mux42 mux42fi34(.a(in34),.b(in70),.c(in106),.d(in142),.sel(cs[1:0]),.out(mux34));
mux42 mux42fi35(.a(in35),.b(in71),.c(in107),.d(in143),.sel(cs[1:0]),.out(mux35));

mux42 mux42fim0(.a(weight0),.b(weight36),.c(weight72),.d(weight108),.sel(cs[1:0]),.out(muxw0));
mux42 mux42fim1(.a(weight1),.b(weight37),.c(weight73),.d(weight109),.sel(cs[1:0]),.out(muxw1));
mux42 mux42fim2(.a(weight2),.b(weight38),.c(weight74),.d(weight110),.sel(cs[1:0]),.out(muxw2));
mux42 mux42fim3(.a(weight3),.b(weight39),.c(weight75),.d(weight111),.sel(cs[1:0]),.out(muxw3));
mux42 mux42fim4(.a(weight4),.b(weight40),.c(weight76),.d(weight112),.sel(cs[1:0]),.out(muxw4));
mux42 mux42fim5(.a(weight5),.b(weight41),.c(weight77),.d(weight113),.sel(cs[1:0]),.out(muxw5));
mux42 mux42fim6(.a(weight6),.b(weight42),.c(weight78),.d(weight114),.sel(cs[1:0]),.out(muxw6));
mux42 mux42fim7(.a(weight7),.b(weight43),.c(weight79),.d(weight115),.sel(cs[1:0]),.out(muxw7));
mux42 mux42fim8(.a(weight8),.b(weight44),.c(weight80),.d(weight116),.sel(cs[1:0]),.out(muxw8));
mux42 mux42fim9(.a(weight9),.b(weight45),.c(weight81),.d(weight117),.sel(cs[1:0]),.out(muxw9));
mux42 mux42fim10(.a(weight10),.b(weight46),.c(weight82),.d(weight118),.sel(cs[1:0]),.out(muxw10));
mux42 mux42fim11(.a(weight11),.b(weight47),.c(weight83),.d(weight119),.sel(cs[1:0]),.out(muxw11));
mux42 mux42fim12(.a(weight12),.b(weight48),.c(weight84),.d(weight120),.sel(cs[1:0]),.out(muxw12));
mux42 mux42fim13(.a(weight13),.b(weight49),.c(weight85),.d(weight121),.sel(cs[1:0]),.out(muxw13));
mux42 mux42fim14(.a(weight14),.b(weight50),.c(weight86),.d(weight122),.sel(cs[1:0]),.out(muxw14));
mux42 mux42fim15(.a(weight15),.b(weight51),.c(weight87),.d(weight123),.sel(cs[1:0]),.out(muxw15));
mux42 mux42fim16(.a(weight16),.b(weight52),.c(weight88),.d(weight124),.sel(cs[1:0]),.out(muxw16));
mux42 mux42fim17(.a(weight17),.b(weight53),.c(weight89),.d(weight125),.sel(cs[1:0]),.out(muxw17));
mux42 mux42fim18(.a(weight18),.b(weight54),.c(weight90),.d(weight126),.sel(cs[1:0]),.out(muxw18));
mux42 mux42fim19(.a(weight19),.b(weight55),.c(weight91),.d(weight127),.sel(cs[1:0]),.out(muxw19));
mux42 mux42fim20(.a(weight20),.b(weight56),.c(weight92),.d(weight128),.sel(cs[1:0]),.out(muxw20));
mux42 mux42fim21(.a(weight21),.b(weight57),.c(weight93),.d(weight129),.sel(cs[1:0]),.out(muxw21));
mux42 mux42fim22(.a(weight22),.b(weight58),.c(weight94),.d(weight130),.sel(cs[1:0]),.out(muxw22));
mux42 mux42fim23(.a(weight23),.b(weight59),.c(weight95),.d(weight131),.sel(cs[1:0]),.out(muxw23));
mux42 mux42fim24(.a(weight24),.b(weight60),.c(weight96),.d(weight132),.sel(cs[1:0]),.out(muxw24));
mux42 mux42fim25(.a(weight25),.b(weight61),.c(weight97),.d(weight133),.sel(cs[1:0]),.out(muxw25));
mux42 mux42fim26(.a(weight26),.b(weight62),.c(weight98),.d(weight134),.sel(cs[1:0]),.out(muxw26));
mux42 mux42fim27(.a(weight27),.b(weight63),.c(weight99),.d(weight135),.sel(cs[1:0]),.out(muxw27));
mux42 mux42fim28(.a(weight28),.b(weight64),.c(weight100),.d(weight136),.sel(cs[1:0]),.out(muxw28));
mux42 mux42fim29(.a(weight29),.b(weight65),.c(weight101),.d(weight137),.sel(cs[1:0]),.out(muxw29));
mux42 mux42fim30(.a(weight30),.b(weight66),.c(weight102),.d(weight138),.sel(cs[1:0]),.out(muxw30));
mux42 mux42fim31(.a(weight31),.b(weight67),.c(weight103),.d(weight139),.sel(cs[1:0]),.out(muxw31));
mux42 mux42fim32(.a(weight32),.b(weight68),.c(weight104),.d(weight140),.sel(cs[1:0]),.out(muxw32));
mux42 mux42fim33(.a(weight33),.b(weight69),.c(weight105),.d(weight141),.sel(cs[1:0]),.out(muxw33));
mux42 mux42fim34(.a(weight34),.b(weight70),.c(weight106),.d(weight142),.sel(cs[1:0]),.out(muxw34));
mux42 mux42fim35(.a(weight35),.b(weight71),.c(weight107),.d(weight143),.sel(cs[1:0]),.out(muxw35));

 multiplier mulf0(.a(mux0),.b(muxw0),.product(mulo0));
multiplier mulf1(.a(mux1),.b(muxw1),.product(mulo1));
multiplier mulf2(.a(mux2),.b(muxw2),.product(mulo2));
multiplier mulf3(.a(mux3),.b(muxw3),.product(mulo3));
multiplier mulf4(.a(mux4),.b(muxw4),.product(mulo4));
multiplier mulf5(.a(mux5),.b(muxw5),.product(mulo5));
multiplier mulf6(.a(mux6),.b(muxw6),.product(mulo6));
multiplier mulf7(.a(mux7),.b(muxw7),.product(mulo7));
multiplier mulf8(.a(mux8),.b(muxw8),.product(mulo8));
multiplier mulf9(.a(mux9),.b(muxw9),.product(mulo9));
multiplier mulf10(.a(mux10),.b(muxw10),.product(mulo10));
multiplier mulf11(.a(mux11),.b(muxw11),.product(mulo11));
multiplier mulf12(.a(mux12),.b(muxw12),.product(mulo12));
multiplier mulf13(.a(mux13),.b(muxw13),.product(mulo13));
multiplier mulf14(.a(mux14),.b(muxw14),.product(mulo14));
multiplier mulf15(.a(mux15),.b(muxw15),.product(mulo15));
multiplier mulf16(.a(mux16),.b(muxw16),.product(mulo16));
multiplier mulf17(.a(mux17),.b(muxw17),.product(mulo17));
multiplier mulf18(.a(mux18),.b(muxw18),.product(mulo18));
multiplier mulf19(.a(mux19),.b(muxw19),.product(mulo19));
multiplier mulf20(.a(mux20),.b(muxw20),.product(mulo20));
multiplier mulf21(.a(mux21),.b(muxw21),.product(mulo21));
multiplier mulf22(.a(mux22),.b(muxw22),.product(mulo22));
multiplier mulf23(.a(mux23),.b(muxw23),.product(mulo23));
multiplier mulf24(.a(mux24),.b(muxw24),.product(mulo24));
multiplier mulf25(.a(mux25),.b(muxw25),.product(mulo25));
multiplier mulf26(.a(mux26),.b(muxw26),.product(mulo26));
multiplier mulf27(.a(mux27),.b(muxw27),.product(mulo27));
multiplier mulf28(.a(mux28),.b(muxw28),.product(mulo28));
multiplier mulf29(.a(mux29),.b(muxw29),.product(mulo29));
multiplier mulf30(.a(mux30),.b(muxw30),.product(mulo30));
multiplier mulf31(.a(mux31),.b(muxw31),.product(mulo31));
multiplier mulf32(.a(mux32),.b(muxw32),.product(mulo32));
multiplier mulf33(.a(mux33),.b(muxw33),.product(mulo33));
multiplier mulf34(.a(mux34),.b(muxw34),.product(mulo34));
multiplier mulf35(.a(mux35),.b(muxw35),.product(mulo35));

/*demux42 demux42fim0(.a(muxo0),.b(muxo36),.c(muxo72),.d(muxo108),.sel(cs[3:2]),.out(mulo0));
demux42 demux42fim1(.a(muxo1),.b(muxo37),.c(muxo73),.d(muxo109),.sel(cs[3:2]),.out(mulo1));
demux42 demux42fim2(.a(muxo2),.b(muxo38),.c(muxo74),.d(muxo110),.sel(cs[3:2]),.out(mulo2));
demux42 demux42fim3(.a(muxo3),.b(muxo39),.c(muxo75),.d(muxo111),.sel(cs[3:2]),.out(mulo3));
demux42 demux42fim4(.a(muxo4),.b(muxo40),.c(muxo76),.d(muxo112),.sel(cs[3:2]),.out(mulo4));
demux42 demux42fim5(.a(muxo5),.b(muxo41),.c(muxo77),.d(muxo113),.sel(cs[3:2]),.out(mulo5));
demux42 demux42fim6(.a(muxo6),.b(muxo42),.c(muxo78),.d(muxo114),.sel(cs[3:2]),.out(mulo6));
demux42 demux42fim7(.a(muxo7),.b(muxo43),.c(muxo79),.d(muxo115),.sel(cs[3:2]),.out(mulo7));
demux42 demux42fim8(.a(muxo8),.b(muxo44),.c(muxo80),.d(muxo116),.sel(cs[3:2]),.out(mulo8));
demux42 demux42fim9(.a(muxo9),.b(muxo45),.c(muxo81),.d(muxo117),.sel(cs[3:2]),.out(mulo9));
demux42 demux42fim10(.a(muxo10),.b(muxo46),.c(muxo82),.d(muxo118),.sel(cs[3:2]),.out(mulo10));
demux42 demux42fim11(.a(muxo11),.b(muxo47),.c(muxo83),.d(muxo119),.sel(cs[3:2]),.out(mulo11));
demux42 demux42fim12(.a(muxo12),.b(muxo48),.c(muxo84),.d(muxo120),.sel(cs[3:2]),.out(mulo12));
demux42 demux42fim13(.a(muxo13),.b(muxo49),.c(muxo85),.d(muxo121),.sel(cs[3:2]),.out(mulo13));
demux42 demux42fim14(.a(muxo14),.b(muxo50),.c(muxo86),.d(muxo122),.sel(cs[3:2]),.out(mulo14));
demux42 demux42fim15(.a(muxo15),.b(muxo51),.c(muxo87),.d(muxo123),.sel(cs[3:2]),.out(mulo15));
demux42 demux42fim16(.a(muxo16),.b(muxo52),.c(muxo88),.d(muxo124),.sel(cs[3:2]),.out(mulo16));
demux42 demux42fim17(.a(muxo17),.b(muxo53),.c(muxo89),.d(muxo125),.sel(cs[3:2]),.out(mulo17));
demux42 demux42fim18(.a(muxo18),.b(muxo54),.c(muxo90),.d(muxo126),.sel(cs[3:2]),.out(mulo18));
demux42 demux42fim19(.a(muxo19),.b(muxo55),.c(muxo91),.d(muxo127),.sel(cs[3:2]),.out(mulo19));
demux42 demux42fim20(.a(muxo20),.b(muxo56),.c(muxo92),.d(muxo128),.sel(cs[3:2]),.out(mulo20));
demux42 demux42fim21(.a(muxo21),.b(muxo57),.c(muxo93),.d(muxo129),.sel(cs[3:2]),.out(mulo21));
demux42 demux42fim22(.a(muxo22),.b(muxo58),.c(muxo94),.d(muxo130),.sel(cs[3:2]),.out(mulo22));
demux42 demux42fim23(.a(muxo23),.b(muxo59),.c(muxo95),.d(muxo131),.sel(cs[3:2]),.out(mulo23));
demux42 demux42fim24(.a(muxo24),.b(muxo60),.c(muxo96),.d(muxo132),.sel(cs[3:2]),.out(mulo24));
demux42 demux42fim25(.a(muxo25),.b(muxo61),.c(muxo97),.d(muxo133),.sel(cs[3:2]),.out(mulo25));
demux42 demux42fim26(.a(muxo26),.b(muxo62),.c(muxo98),.d(muxo134),.sel(cs[3:2]),.out(mulo26));
demux42 demux42fim27(.a(muxo27),.b(muxo63),.c(muxo99),.d(muxo135),.sel(cs[3:2]),.out(mulo27));
demux42 demux42fim28(.a(muxo28),.b(muxo64),.c(muxo100),.d(muxo136),.sel(cs[3:2]),.out(mulo28));
demux42 demux42fim29(.a(muxo29),.b(muxo65),.c(muxo101),.d(muxo137),.sel(cs[3:2]),.out(mulo29));
demux42 demux42fim30(.a(muxo30),.b(muxo66),.c(muxo102),.d(muxo138),.sel(cs[3:2]),.out(mulo30));
demux42 demux42fim31(.a(muxo31),.b(muxo67),.c(muxo103),.d(muxo139),.sel(cs[3:2]),.out(mulo31));
demux42 demux42fim32(.a(muxo32),.b(muxo68),.c(muxo104),.d(muxo140),.sel(cs[3:2]),.out(mulo32));
demux42 demux42fim33(.a(muxo33),.b(muxo69),.c(muxo105),.d(muxo141),.sel(cs[3:2]),.out(mulo33));
demux42 demux42fim34(.a(muxo34),.b(muxo70),.c(muxo106),.d(muxo142),.sel(cs[3:2]),.out(mulo34));
demux42 demux42fim35(.a(muxo35),.b(muxo71),.c(muxo107),.d(muxo143),.sel(cs[3:2]),.out(mulo35));
*/
reg [7:0] mulreg0;
reg [7:0] mulreg1;
reg [7:0] mulreg2;
reg [7:0] mulreg3;
reg [7:0] mulreg4;
reg [7:0] mulreg5;
reg [7:0] mulreg6;
reg [7:0] mulreg7;
reg [7:0] mulreg8;
reg [7:0] mulreg9;
reg [7:0] mulreg10;
reg [7:0] mulreg11;
reg [7:0] mulreg12;
reg [7:0] mulreg13;
reg [7:0] mulreg14;
reg [7:0] mulreg15;
reg [7:0] mulreg16;
reg [7:0] mulreg17;
reg [7:0] mulreg18;
reg [7:0] mulreg19;
reg [7:0] mulreg20;
reg [7:0] mulreg21;
reg [7:0] mulreg22;
reg [7:0] mulreg23;
reg [7:0] mulreg24;
reg [7:0] mulreg25;
reg [7:0] mulreg26;
reg [7:0] mulreg27;
reg [7:0] mulreg28;
reg [7:0] mulreg29;
reg [7:0] mulreg30;
reg [7:0] mulreg31;
reg [7:0] mulreg32;
reg [7:0] mulreg33;
reg [7:0] mulreg34;
reg [7:0] mulreg35;
reg [7:0] mulreg36;
reg [7:0] mulreg37;
reg [7:0] mulreg38;
reg [7:0] mulreg39;
reg [7:0] mulreg40;
reg [7:0] mulreg41;
reg [7:0] mulreg42;
reg [7:0] mulreg43;
reg [7:0] mulreg44;
reg [7:0] mulreg45;
reg [7:0] mulreg46;
reg [7:0] mulreg47;
reg [7:0] mulreg48;
reg [7:0] mulreg49;
reg [7:0] mulreg50;
reg [7:0] mulreg51;
reg [7:0] mulreg52;
reg [7:0] mulreg53;
reg [7:0] mulreg54;
reg [7:0] mulreg55;
reg [7:0] mulreg56;
reg [7:0] mulreg57;
reg [7:0] mulreg58;
reg [7:0] mulreg59;
reg [7:0] mulreg60;
reg [7:0] mulreg61;
reg [7:0] mulreg62;
reg [7:0] mulreg63;
reg [7:0] mulreg64;
reg [7:0] mulreg65;
reg [7:0] mulreg66;
reg [7:0] mulreg67;
reg [7:0] mulreg68;
reg [7:0] mulreg69;
reg [7:0] mulreg70;
reg [7:0] mulreg71;
reg [7:0] mulreg72;
reg [7:0] mulreg73;
reg [7:0] mulreg74;
reg [7:0] mulreg75;
reg [7:0] mulreg76;
reg [7:0] mulreg77;
reg [7:0] mulreg78;
reg [7:0] mulreg79;
reg [7:0] mulreg80;
reg [7:0] mulreg81;
reg [7:0] mulreg82;
reg [7:0] mulreg83;
reg [7:0] mulreg84;
reg [7:0] mulreg85;
reg [7:0] mulreg86;
reg [7:0] mulreg87;
reg [7:0] mulreg88;
reg [7:0] mulreg89;
reg [7:0] mulreg90;
reg [7:0] mulreg91;
reg [7:0] mulreg92;
reg [7:0] mulreg93;
reg [7:0] mulreg94;
reg [7:0] mulreg95;
reg [7:0] mulreg96;
reg [7:0] mulreg97;
reg [7:0] mulreg98;
reg [7:0] mulreg99;
reg [7:0] mulreg100;
reg [7:0] mulreg101;
reg [7:0] mulreg102;
reg [7:0] mulreg103;
reg [7:0] mulreg104;
reg [7:0] mulreg105;
reg [7:0] mulreg106;
reg [7:0] mulreg107;
reg [7:0] mulreg108;
reg [7:0] mulreg109;
reg [7:0] mulreg110;
reg [7:0] mulreg111;
reg [7:0] mulreg112;
reg [7:0] mulreg113;
reg [7:0] mulreg114;
reg [7:0] mulreg115;
reg [7:0] mulreg116;
reg [7:0] mulreg117;
reg [7:0] mulreg118;
reg [7:0] mulreg119;
reg [7:0] mulreg120;
reg [7:0] mulreg121;
reg [7:0] mulreg122;
reg [7:0] mulreg123;
reg [7:0] mulreg124;
reg [7:0] mulreg125;
reg [7:0] mulreg126;
reg [7:0] mulreg127;
reg [7:0] mulreg128;
reg [7:0] mulreg129;
reg [7:0] mulreg130;
reg [7:0] mulreg131;
reg [7:0] mulreg132;
reg [7:0] mulreg133;
reg [7:0] mulreg134;
reg [7:0] mulreg135;
reg [7:0] mulreg136;
reg [7:0] mulreg137;
reg [7:0] mulreg138;
reg [7:0] mulreg139;
reg [7:0] mulreg140;
reg [7:0] mulreg141;
reg [7:0] mulreg142;
reg [7:0] mulreg143;

 
reg [7:0] outreg;

wire [7:0] outadd1; 

reg [2:0] state;
localparam WAIT = 3'b000;
localparam CALCM1 = 3'b001;
localparam CALCM2 = 3'b010;
localparam CALCM3 = 3'b011;
localparam CALCM4 = 3'b100;
localparam CALC2  = 3'b101;
localparam READY = 3'b110;
localparam START = 3'b111;
reg [2:0] next_state;


adderF adderf1(.in0(mulreg0),.in1(mulreg1),.in2(mulreg2),.in3(mulreg3),.in4(mulreg4),.in5(mulreg5),.in6(mulreg6),.in7(mulreg7),.in8(mulreg8),.in9(mulreg9),.in10(mulreg10),.in11(mulreg11),.in12(mulreg12),.in13(mulreg13),.in14(mulreg14),.in15(mulreg15),.in16(mulreg16),.in17(mulreg17),.in18(mulreg18),.in19(mulreg19),.in20(mulreg20),.in21(mulreg21),.in22(mulreg22),.in23(mulreg23),.in24(mulreg24),.in25(mulreg25),.in26(mulreg26),.in27(mulreg27),.in28(mulreg28),.in29(mulreg29),.in30(mulreg30),.in31(mulreg31),.in32(mulreg32),.in33(mulreg33),.in34(mulreg34),.in35(mulreg35),.in36(mulreg36),.in37(mulreg37),.in38(mulreg38),.in39(mulreg39),.in40(mulreg40),.in41(mulreg41),.in42(mulreg42),.in43(mulreg43),.in44(mulreg44),.in45(mulreg45),.in46(mulreg46),.in47(mulreg47),.in48(mulreg48),.in49(mulreg49),.in50(mulreg50),.in51(mulreg51),.in52(mulreg52),.in53(mulreg53),.in54(mulreg54),.in55(mulreg55),.in56(mulreg56),.in57(mulreg57),.in58(mulreg58),.in59(mulreg59),.in60(mulreg60),.in61(mulreg61),.in62(mulreg62),.in63(mulreg63),.in64(mulreg64),.in65(mulreg65),.in66(mulreg66),.in67(mulreg67),.in68(mulreg68),.in69(mulreg69),.in70(mulreg70),.in71(mulreg71),.in72(mulreg72),.in73(mulreg73),.in74(mulreg74),.in75(mulreg75),.in76(mulreg76),.in77(mulreg77),.in78(mulreg78),.in79(mulreg79),.in80(mulreg80),.in81(mulreg81),.in82(mulreg82),.in83(mulreg83),.in84(mulreg84),.in85(mulreg85),.in86(mulreg86),.in87(mulreg87),.in88(mulreg88),.in89(mulreg89),.in90(mulreg90),.in91(mulreg91),.in92(mulreg92),.in93(mulreg93),.in94(mulreg94),.in95(mulreg95),.in96(mulreg96),.in97(mulreg97),.in98(mulreg98),.in99(mulreg99),.in100(mulreg100),.in101(mulreg101),.in102(mulreg102),.in103(mulreg103),.in104(mulreg104),.in105(mulreg105),.in106(mulreg106),.in107(mulreg107),.in108(mulreg108),.in109(mulreg109),.in110(mulreg110),.in111(mulreg111),.in112(mulreg112),.in113(mulreg113),.in114(mulreg114),.in115(mulreg115),.in116(mulreg116),.in117(mulreg117),.in118(mulreg118),.in119(mulreg119),.in120(mulreg120),.in121(mulreg121),.in122(mulreg122),.in123(mulreg123),.in124(mulreg124),.in125(mulreg125),.in126(mulreg126),.in127(mulreg127),.in128(mulreg128),.in129(mulreg129),.in130(mulreg130),.in131(mulreg131),.in132(mulreg132),.in133(mulreg133),.in134(mulreg134),.in135(mulreg135),.in136(mulreg136),.in137(mulreg137),.in138(mulreg138),.in139(mulreg139),.in140(mulreg140),.in141(mulreg141),.in142(mulreg142),.in143(mulreg143),
.out(outadd1));

always @(posedge clk or posedge start)
begin
	if (start) begin
	$monitor("%b",state);
	next_state <= START;
	ready <= 0;
	end
	else state <= next_state;
	case (state)
		START:
		begin 
		next_state <= CALCM1;
		cs <= 4'b0000;
		ready <= 0;
		end
		CALCM1:
		begin 
		mulreg0<=mulo0;mulreg1<=mulo1;mulreg2<=mulo2;mulreg3<=mulo3;mulreg4<=mulo4;mulreg5<=mulo5;mulreg6<=mulo6;mulreg7<=mulo7;mulreg8<=mulo8;mulreg9<=mulo9;mulreg10<=mulo10;mulreg11<=mulo11;mulreg12<=mulo12;mulreg13<=mulo13;mulreg14<=mulo14;mulreg15<=mulo15;mulreg16<=mulo16;mulreg17<=mulo17;mulreg18<=mulo18;mulreg19<=mulo19;mulreg20<=mulo20;mulreg21<=mulo21;mulreg22<=mulo22;mulreg23<=mulo23;mulreg24<=mulo24;mulreg25<=mulo25;mulreg26<=mulo26;mulreg27<=mulo27;mulreg28<=mulo28;mulreg29<=mulo29;mulreg30<=mulo30;mulreg31<=mulo31;mulreg32<=mulo32;mulreg33<=mulo33;mulreg34<=mulo34;mulreg35<=mulo35;
		next_state <= CALCM2;
		cs <= 4'b0101;
		end
		CALCM2:
		begin 
		next_state <= CALCM3;
		mulreg36<=mulo0;mulreg37<=mulo1;mulreg38<=mulo2;mulreg39<=mulo3;mulreg40<=mulo4;mulreg41<=mulo5;mulreg42<=mulo6;mulreg43<=mulo7;mulreg44<=mulo8;mulreg45<=mulo9;mulreg46<=mulo10;mulreg47<=mulo11;mulreg48<=mulo12;mulreg49<=mulo13;mulreg50<=mulo14;mulreg51<=mulo15;mulreg52<=mulo16;mulreg53<=mulo17;mulreg54<=mulo18;mulreg55<=mulo19;mulreg56<=mulo20;mulreg57<=mulo21;mulreg58<=mulo22;mulreg59<=mulo23;mulreg60<=mulo24;mulreg61<=mulo25;mulreg62<=mulo26;mulreg63<=mulo27;mulreg64<=mulo28;mulreg65<=mulo29;mulreg66<=mulo30;mulreg67<=mulo31;mulreg68<=mulo32;mulreg69<=mulo33;mulreg70<=mulo34;mulreg71<=mulo35;
		cs <= 4'b1010;
		end
		CALCM3:
		begin 
		next_state <= CALCM4;
		mulreg72<=mulo0;mulreg73<=mulo1;mulreg74<=mulo2;mulreg75<=mulo3;mulreg76<=mulo4;mulreg77<=mulo5;mulreg78<=mulo6;mulreg79<=mulo7;mulreg80<=mulo8;mulreg81<=mulo9;mulreg82<=mulo10;mulreg83<=mulo11;mulreg84<=mulo12;mulreg85<=mulo13;mulreg86<=mulo14;mulreg87<=mulo15;mulreg88<=mulo16;mulreg89<=mulo17;mulreg90<=mulo18;mulreg91<=mulo19;mulreg92<=mulo20;mulreg93<=mulo21;mulreg94<=mulo22;mulreg95<=mulo23;mulreg96<=mulo24;mulreg97<=mulo25;mulreg98<=mulo26;mulreg99<=mulo27;mulreg100<=mulo28;mulreg101<=mulo29;mulreg102<=mulo30;mulreg103<=mulo31;mulreg104<=mulo32;mulreg105<=mulo33;mulreg106<=mulo34;mulreg107<=mulo35;
		cs <= 4'b1111;
		end
		CALCM4:
		begin 
		next_state <= CALC2;
		mulreg108<=mulo0;mulreg109<=mulo1;mulreg110<=mulo2;mulreg111<=mulo3;mulreg112<=mulo4;mulreg113<=mulo5;mulreg114<=mulo6;mulreg115<=mulo7;mulreg116<=mulo8;mulreg117<=mulo9;mulreg118<=mulo10;mulreg119<=mulo11;mulreg120<=mulo12;mulreg121<=mulo13;mulreg122<=mulo14;mulreg123<=mulo15;mulreg124<=mulo16;mulreg125<=mulo17;mulreg126<=mulo18;mulreg127<=mulo19;mulreg128<=mulo20;mulreg129<=mulo21;mulreg130<=mulo22;mulreg131<=mulo23;mulreg132<=mulo24;mulreg133<=mulo25;mulreg134<=mulo26;mulreg135<=mulo27;mulreg136<=mulo28;mulreg137<=mulo29;mulreg138<=mulo30;mulreg139<=mulo31;mulreg140<=mulo32;mulreg141<=mulo33;mulreg142<=mulo34;mulreg143<=mulo35;
		cs <= 4'b0000;
		end
		CALC2:
		begin 
		next_state <= READY;
		outreg <= outadd1;
		cs <= 4'b0000;
		ready <= 1;
		end
		READY:
		begin 
		next_state <= WAIT;
		cs <= 4'b0000;
		ready <= 0;
		end
		/*default:
		begin 
		state <= WAIT;
		cs <= 4'b0000;
		end*/
	endcase
end 

endmodule

module  adderF(in0,in1,in2,in3,in4,in5,in6,in7,in8,in9,in10,in11,in12,in13,in14,in15,in16,in17,in18,in19,in20,in21,in22,in23,in24,in25,in26,in27,in28,in29,in30,in31,in32,in33,in34,in35,in36,in37,in38,in39,in40,in41,in42,in43,in44,in45,in46,in47,in48,in49,in50,in51,in52,in53,in54,in55,in56,in57,in58,in59,in60,in61,in62,in63,in64,in65,in66,in67,in68,in69,in70,in71,in72,in73,in74,in75,in76,in77,in78,in79,in80,in81,in82,in83,in84,in85,in86,in87,in88,in89,in90,in91,in92,in93,in94,in95,in96,in97,in98,in99,in100,in101,in102,in103,in104,in105,in106,in107,in108,in109,in110,in111,in112,in113,in114,in115,in116,in117,in118,in119,in120,in121,in122,in123,in124,in125,in126,in127,in128,in129,in130,in131,in132,in133,in134,in135,in136,in137,in138,in139,in140,in141,in142,in143,
out);

input [7:0] in0;
input [7:0] in1;
input [7:0] in2;
input [7:0] in3;
input [7:0] in4;
input [7:0] in5;
input [7:0] in6;
input [7:0] in7;
input [7:0] in8;
input [7:0] in9;
input [7:0] in10;
input [7:0] in11;
input [7:0] in12;
input [7:0] in13;
input [7:0] in14;
input [7:0] in15;
input [7:0] in16;
input [7:0] in17;
input [7:0] in18;
input [7:0] in19;
input [7:0] in20;
input [7:0] in21;
input [7:0] in22;
input [7:0] in23;
input [7:0] in24;
input [7:0] in25;
input [7:0] in26;
input [7:0] in27;
input [7:0] in28;
input [7:0] in29;
input [7:0] in30;
input [7:0] in31;
input [7:0] in32;
input [7:0] in33;
input [7:0] in34;
input [7:0] in35;
input [7:0] in36;
input [7:0] in37;
input [7:0] in38;
input [7:0] in39;
input [7:0] in40;
input [7:0] in41;
input [7:0] in42;
input [7:0] in43;
input [7:0] in44;
input [7:0] in45;
input [7:0] in46;
input [7:0] in47;
input [7:0] in48;
input [7:0] in49;
input [7:0] in50;
input [7:0] in51;
input [7:0] in52;
input [7:0] in53;
input [7:0] in54;
input [7:0] in55;
input [7:0] in56;
input [7:0] in57;
input [7:0] in58;
input [7:0] in59;
input [7:0] in60;
input [7:0] in61;
input [7:0] in62;
input [7:0] in63;
input [7:0] in64;
input [7:0] in65;
input [7:0] in66;
input [7:0] in67;
input [7:0] in68;
input [7:0] in69;
input [7:0] in70;
input [7:0] in71;
input [7:0] in72;
input [7:0] in73;
input [7:0] in74;
input [7:0] in75;
input [7:0] in76;
input [7:0] in77;
input [7:0] in78;
input [7:0] in79;
input [7:0] in80;
input [7:0] in81;
input [7:0] in82;
input [7:0] in83;
input [7:0] in84;
input [7:0] in85;
input [7:0] in86;
input [7:0] in87;
input [7:0] in88;
input [7:0] in89;
input [7:0] in90;
input [7:0] in91;
input [7:0] in92;
input [7:0] in93;
input [7:0] in94;
input [7:0] in95;
input [7:0] in96;
input [7:0] in97;
input [7:0] in98;
input [7:0] in99;
input [7:0] in100;
input [7:0] in101;
input [7:0] in102;
input [7:0] in103;
input [7:0] in104;
input [7:0] in105;
input [7:0] in106;
input [7:0] in107;
input [7:0] in108;
input [7:0] in109;
input [7:0] in110;
input [7:0] in111;
input [7:0] in112;
input [7:0] in113;
input [7:0] in114;
input [7:0] in115;
input [7:0] in116;
input [7:0] in117;
input [7:0] in118;
input [7:0] in119;
input [7:0] in120;
input [7:0] in121;
input [7:0] in122;
input [7:0] in123;
input [7:0] in124;
input [7:0] in125;
input [7:0] in126;
input [7:0] in127;
input [7:0] in128;
input [7:0] in129;
input [7:0] in130;
input [7:0] in131;
input [7:0] in132;
input [7:0] in133;
input [7:0] in134;
input [7:0] in135;
input [7:0] in136;
input [7:0] in137;
input [7:0] in138;
input [7:0] in139;
input [7:0] in140;
input [7:0] in141;
input [7:0] in142;
input [7:0] in143;
output [7:0] out;

assign out =  in0+in1+in2+in3+in4+in5+in6+in7+in8+in9+in10+in11+in12+in13+in14+in15+in16+in17+in18+in19+in20+in21+in22+in23+in24+in25+in26+in27+in28+in29+in30+in31+in32+in33+in34+in35+in36+in37+in38+in39+in40+in41+in42+in43+in44+in45+in46+in47+in48+in49+in50+in51+in52+in53+in54+in55+in56+in57+in58+in59+in60+in61+in62+in63+in64+in65+in66+in67+in68+in69+in70+in71+in72+in73+in74+in75+in76+in77+in78+in79+in80+in81+in82+in83+in84+in85+in86+in87+in88+in89+in90+in91+in92+in93+in94+in95+in96+in97+in98+in99+in100+in101+in102+in103+in104+in105+in106+in107+in108+in109+in110+in111+in112+in113+in114+in115+in116+in117+in118+in119+in120+in121+in122+in123+in124+in125+in126+in127+in128+in129+in130+in131+in132+in133+in134+in135+in136+in137+in138+in139+in140+in141+in142+in143;

endmodule