`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    13:15:54 11/05/2017 
// Design Name: 
// Module Name:    poolinglayer 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module poolinglayer( in0,in1,in2,in3,in4,in5,in6,in7,in8,in9,in10,in11,in12,in13,in14,
in15,in16,in17,in18,in19,in20,in21,in22,in23,in24,in25,in26,in27,in28,in29,in30,in31,
in32,in33,in34,in35,in36,in37,in38,in39,in40,in41,in42,in43,in44,in45,in46,in47,in48,
in49,in50,in51,in52,in53,in54,in55,in56,in57,in58,in59,in60,in61,in62,in63,in64,in65,
in66,in67,in68,in69,in70,in71,in72,in73,in74,in75,in76,in77,in78,in79,in80,in81,in82,
in83,in84,in85,in86,in87,in88,in89,in90,in91,in92,in93,in94,in95,in96,in97,in98,in99,
in100,in101,in102,in103,in104,in105,in106,in107,in108,in109,in110,in111,in112,in113,
in114,in115,in116,in117,in118,in119,in120,in121,in122,in123,in124,in125,in126,in127,
in128,in129,in130,in131,in132,in133,in134,in135,in136,in137,in138,in139,in140,in141,
in142,in143,in144,in145,in146,in147,in148,in149,in150,in151,in152,in153,in154,in155,
in156,in157,in158,in159,in160,in161,in162,in163,in164,in165,in166,in167,in168,in169,
in170,in171,in172,in173,in174,in175,in176,in177,in178,in179,in180,in181,in182,in183,
in184,in185,in186,in187,in188,in189,in190,in191,in192,in193,in194,in195,in196,in197,
in198,in199,in200,in201,in202,in203,in204,in205,in206,in207,in208,in209,in210,in211,
in212,in213,in214,in215,in216,in217,in218,in219,in220,in221,in222,in223,in224,in225,
in226,in227,in228,in229,in230,in231,in232,in233,in234,in235,in236,in237,in238,in239,
in240,in241,in242,in243,in244,in245,in246,in247,in248,in249,in250,in251,in252,in253,
in254,in255,in256,in257,in258,in259,in260,in261,in262,in263,in264,in265,in266,in267,
in268,in269,in270,in271,in272,in273,in274,in275,in276,in277,in278,in279,in280,in281,
in282,in283,in284,in285,in286,in287,in288,in289,in290,in291,in292,in293,in294,in295,
in296,in297,in298,in299,in300,in301,in302,in303,in304,in305,in306,in307,in308,in309,
in310,in311,in312,in313,in314,in315,in316,in317,in318,in319,in320,in321,in322,in323,
in324,in325,in326,in327,in328,in329,in330,in331,in332,in333,in334,in335,in336,in337,
in338,in339,in340,in341,in342,in343,in344,in345,in346,in347,in348,in349,in350,in351,in352,
in353,in354,in355,in356,in357,in358,in359,in360,in361,in362,in363,in364,in365,in366,
in367,in368,in369,in370,in371,in372,in373,in374,in375,in376,in377,in378,in379,in380,
in381,in382,in383,in384,in385,in386,in387,in388,in389,in390,in391,in392,in393,in394,
in395,in396,in397,in398,in399,in400,in401,in402,in403,in404,in405,in406,in407,in408,
in409,in410,in411,in412,in413,in414,in415,in416,in417,in418,in419,in420,in421,in422,
in423,in424,in425,in426,in427,in428,in429,in430,in431,in432,in433,in434,in435,in436,
in437,in438,in439,in440,in441,in442,in443,in444,in445,in446,in447,in448,in449,in450,
in451,in452,in453,in454,in455,in456,in457,in458,in459,in460,in461,in462,in463,in464,
in465,in466,in467,in468,in469,in470,in471,in472,in473,in474,in475,in476,in477,in478,
in479,in480,in481,in482,in483,in484,in485,in486,in487,in488,in489,in490,in491,in492,
in493,in494,in495,in496,in497,in498,in499,in500,in501,in502,in503,in504,in505,in506,
in507,in508,in509,in510,in511,in512,in513,in514,in515,in516,in517,in518,in519,in520,
in521,in522,in523,in524,in525,in526,in527,in528,in529,in530,in531,in532,in533,in534,
in535,in536,in537,in538,in539,in540,in541,in542,in543,in544,in545,in546,in547,in548,
in549,in550,in551,in552,in553,in554,in555,in556,in557,in558,in559,in560,in561,in562,
in563,in564,in565,in566,in567,in568,in569,in570,in571,in572,in573,in574,in575, out0,out1,out2,out3,out4,out5,out6,out7,out8,out9,out10,out11,out12,out13,out14,out15,out16,out17,out18,out19,out20,out21,out22,out23,out24,out25,out26,out27,out28,out29,out30,out31,out32,out33,out34,out35,out36,out37,out38,out39,out40,out41,out42,out43,out44,out45,out46,out47,out48,out49,out50,out51,out52,out53,out54,out55,out56,out57,out58,out59,out60,out61,out62,out63,out64,out65,out66,out67,out68,out69,out70,out71,out72,out73,out74,out75,out76,out77,out78,out79,out80,out81,out82,out83,out84,out85,out86,out87,out88,out89,out90,out91,out92,out93,out94,out95,out96,out97,out98,out99,out100,out101,out102,out103,out104,out105,out106,out107,out108,out109,out110,out111,out112,out113,out114,out115,out116,out117,out118,out119,out120,out121,out122,out123,out124,out125,out126,out127,out128,out129,out130,out131,out132,out133,out134,out135,out136,out137,out138,out139,out140,out141,out142,out143
,clk,ready,start);

input clk;
input start;
 input [7:0] in0;
input [7:0] in1;
input [7:0] in2;
input [7:0] in3;
input [7:0] in4;
input [7:0] in5;
input [7:0] in6;
input [7:0] in7;
input [7:0] in8;
input [7:0] in9;
input [7:0] in10;
input [7:0] in11;
input [7:0] in12;
input [7:0] in13;
input [7:0] in14;
input [7:0] in15;
input [7:0] in16;
input [7:0] in17;
input [7:0] in18;
input [7:0] in19;
input [7:0] in20;
input [7:0] in21;
input [7:0] in22;
input [7:0] in23;
input [7:0] in24;
input [7:0] in25;
input [7:0] in26;
input [7:0] in27;
input [7:0] in28;
input [7:0] in29;
input [7:0] in30;
input [7:0] in31;
input [7:0] in32;
input [7:0] in33;
input [7:0] in34;
input [7:0] in35;
input [7:0] in36;
input [7:0] in37;
input [7:0] in38;
input [7:0] in39;
input [7:0] in40;
input [7:0] in41;
input [7:0] in42;
input [7:0] in43;
input [7:0] in44;
input [7:0] in45;
input [7:0] in46;
input [7:0] in47;
input [7:0] in48;
input [7:0] in49;
input [7:0] in50;
input [7:0] in51;
input [7:0] in52;
input [7:0] in53;
input [7:0] in54;
input [7:0] in55;
input [7:0] in56;
input [7:0] in57;
input [7:0] in58;
input [7:0] in59;
input [7:0] in60;
input [7:0] in61;
input [7:0] in62;
input [7:0] in63;
input [7:0] in64;
input [7:0] in65;
input [7:0] in66;
input [7:0] in67;
input [7:0] in68;
input [7:0] in69;
input [7:0] in70;
input [7:0] in71;
input [7:0] in72;
input [7:0] in73;
input [7:0] in74;
input [7:0] in75;
input [7:0] in76;
input [7:0] in77;
input [7:0] in78;
input [7:0] in79;
input [7:0] in80;
input [7:0] in81;
input [7:0] in82;
input [7:0] in83;
input [7:0] in84;
input [7:0] in85;
input [7:0] in86;
input [7:0] in87;
input [7:0] in88;
input [7:0] in89;
input [7:0] in90;
input [7:0] in91;
input [7:0] in92;
input [7:0] in93;
input [7:0] in94;
input [7:0] in95;
input [7:0] in96;
input [7:0] in97;
input [7:0] in98;
input [7:0] in99;
input [7:0] in100;
input [7:0] in101;
input [7:0] in102;
input [7:0] in103;
input [7:0] in104;
input [7:0] in105;
input [7:0] in106;
input [7:0] in107;
input [7:0] in108;
input [7:0] in109;
input [7:0] in110;
input [7:0] in111;
input [7:0] in112;
input [7:0] in113;
input [7:0] in114;
input [7:0] in115;
input [7:0] in116;
input [7:0] in117;
input [7:0] in118;
input [7:0] in119;
input [7:0] in120;
input [7:0] in121;
input [7:0] in122;
input [7:0] in123;
input [7:0] in124;
input [7:0] in125;
input [7:0] in126;
input [7:0] in127;
input [7:0] in128;
input [7:0] in129;
input [7:0] in130;
input [7:0] in131;
input [7:0] in132;
input [7:0] in133;
input [7:0] in134;
input [7:0] in135;
input [7:0] in136;
input [7:0] in137;
input [7:0] in138;
input [7:0] in139;
input [7:0] in140;
input [7:0] in141;
input [7:0] in142;
input [7:0] in143;
input [7:0] in144;
input [7:0] in145;
input [7:0] in146;
input [7:0] in147;
input [7:0] in148;
input [7:0] in149;
input [7:0] in150;
input [7:0] in151;
input [7:0] in152;
input [7:0] in153;
input [7:0] in154;
input [7:0] in155;
input [7:0] in156;
input [7:0] in157;
input [7:0] in158;
input [7:0] in159;
input [7:0] in160;
input [7:0] in161;
input [7:0] in162;
input [7:0] in163;
input [7:0] in164;
input [7:0] in165;
input [7:0] in166;
input [7:0] in167;
input [7:0] in168;
input [7:0] in169;
input [7:0] in170;
input [7:0] in171;
input [7:0] in172;
input [7:0] in173;
input [7:0] in174;
input [7:0] in175;
input [7:0] in176;
input [7:0] in177;
input [7:0] in178;
input [7:0] in179;
input [7:0] in180;
input [7:0] in181;
input [7:0] in182;
input [7:0] in183;
input [7:0] in184;
input [7:0] in185;
input [7:0] in186;
input [7:0] in187;
input [7:0] in188;
input [7:0] in189;
input [7:0] in190;
input [7:0] in191;
input [7:0] in192;
input [7:0] in193;
input [7:0] in194;
input [7:0] in195;
input [7:0] in196;
input [7:0] in197;
input [7:0] in198;
input [7:0] in199;
input [7:0] in200;
input [7:0] in201;
input [7:0] in202;
input [7:0] in203;
input [7:0] in204;
input [7:0] in205;
input [7:0] in206;
input [7:0] in207;
input [7:0] in208;
input [7:0] in209;
input [7:0] in210;
input [7:0] in211;
input [7:0] in212;
input [7:0] in213;
input [7:0] in214;
input [7:0] in215;
input [7:0] in216;
input [7:0] in217;
input [7:0] in218;
input [7:0] in219;
input [7:0] in220;
input [7:0] in221;
input [7:0] in222;
input [7:0] in223;
input [7:0] in224;
input [7:0] in225;
input [7:0] in226;
input [7:0] in227;
input [7:0] in228;
input [7:0] in229;
input [7:0] in230;
input [7:0] in231;
input [7:0] in232;
input [7:0] in233;
input [7:0] in234;
input [7:0] in235;
input [7:0] in236;
input [7:0] in237;
input [7:0] in238;
input [7:0] in239;
input [7:0] in240;
input [7:0] in241;
input [7:0] in242;
input [7:0] in243;
input [7:0] in244;
input [7:0] in245;
input [7:0] in246;
input [7:0] in247;
input [7:0] in248;
input [7:0] in249;
input [7:0] in250;
input [7:0] in251;
input [7:0] in252;
input [7:0] in253;
input [7:0] in254;
input [7:0] in255;
input [7:0] in256;
input [7:0] in257;
input [7:0] in258;
input [7:0] in259;
input [7:0] in260;
input [7:0] in261;
input [7:0] in262;
input [7:0] in263;
input [7:0] in264;
input [7:0] in265;
input [7:0] in266;
input [7:0] in267;
input [7:0] in268;
input [7:0] in269;
input [7:0] in270;
input [7:0] in271;
input [7:0] in272;
input [7:0] in273;
input [7:0] in274;
input [7:0] in275;
input [7:0] in276;
input [7:0] in277;
input [7:0] in278;
input [7:0] in279;
input [7:0] in280;
input [7:0] in281;
input [7:0] in282;
input [7:0] in283;
input [7:0] in284;
input [7:0] in285;
input [7:0] in286;
input [7:0] in287;
input [7:0] in288;
input [7:0] in289;
input [7:0] in290;
input [7:0] in291;
input [7:0] in292;
input [7:0] in293;
input [7:0] in294;
input [7:0] in295;
input [7:0] in296;
input [7:0] in297;
input [7:0] in298;
input [7:0] in299;
input [7:0] in300;
input [7:0] in301;
input [7:0] in302;
input [7:0] in303;
input [7:0] in304;
input [7:0] in305;
input [7:0] in306;
input [7:0] in307;
input [7:0] in308;
input [7:0] in309;
input [7:0] in310;
input [7:0] in311;
input [7:0] in312;
input [7:0] in313;
input [7:0] in314;
input [7:0] in315;
input [7:0] in316;
input [7:0] in317;
input [7:0] in318;
input [7:0] in319;
input [7:0] in320;
input [7:0] in321;
input [7:0] in322;
input [7:0] in323;
input [7:0] in324;
input [7:0] in325;
input [7:0] in326;
input [7:0] in327;
input [7:0] in328;
input [7:0] in329;
input [7:0] in330;
input [7:0] in331;
input [7:0] in332;
input [7:0] in333;
input [7:0] in334;
input [7:0] in335;
input [7:0] in336;
input [7:0] in337;
input [7:0] in338;
input [7:0] in339;
input [7:0] in340;
input [7:0] in341;
input [7:0] in342;
input [7:0] in343;
input [7:0] in344;
input [7:0] in345;
input [7:0] in346;
input [7:0] in347;
input [7:0] in348;
input [7:0] in349;
input [7:0] in350;
input [7:0] in351;
input [7:0] in352;
input [7:0] in353;
input [7:0] in354;
input [7:0] in355;
input [7:0] in356;
input [7:0] in357;
input [7:0] in358;
input [7:0] in359;
input [7:0] in360;
input [7:0] in361;
input [7:0] in362;
input [7:0] in363;
input [7:0] in364;
input [7:0] in365;
input [7:0] in366;
input [7:0] in367;
input [7:0] in368;
input [7:0] in369;
input [7:0] in370;
input [7:0] in371;
input [7:0] in372;
input [7:0] in373;
input [7:0] in374;
input [7:0] in375;
input [7:0] in376;
input [7:0] in377;
input [7:0] in378;
input [7:0] in379;
input [7:0] in380;
input [7:0] in381;
input [7:0] in382;
input [7:0] in383;
input [7:0] in384;
input [7:0] in385;
input [7:0] in386;
input [7:0] in387;
input [7:0] in388;
input [7:0] in389;
input [7:0] in390;
input [7:0] in391;
input [7:0] in392;
input [7:0] in393;
input [7:0] in394;
input [7:0] in395;
input [7:0] in396;
input [7:0] in397;
input [7:0] in398;
input [7:0] in399;
input [7:0] in400;
input [7:0] in401;
input [7:0] in402;
input [7:0] in403;
input [7:0] in404;
input [7:0] in405;
input [7:0] in406;
input [7:0] in407;
input [7:0] in408;
input [7:0] in409;
input [7:0] in410;
input [7:0] in411;
input [7:0] in412;
input [7:0] in413;
input [7:0] in414;
input [7:0] in415;
input [7:0] in416;
input [7:0] in417;
input [7:0] in418;
input [7:0] in419;
input [7:0] in420;
input [7:0] in421;
input [7:0] in422;
input [7:0] in423;
input [7:0] in424;
input [7:0] in425;
input [7:0] in426;
input [7:0] in427;
input [7:0] in428;
input [7:0] in429;
input [7:0] in430;
input [7:0] in431;
input [7:0] in432;
input [7:0] in433;
input [7:0] in434;
input [7:0] in435;
input [7:0] in436;
input [7:0] in437;
input [7:0] in438;
input [7:0] in439;
input [7:0] in440;
input [7:0] in441;
input [7:0] in442;
input [7:0] in443;
input [7:0] in444;
input [7:0] in445;
input [7:0] in446;
input [7:0] in447;
input [7:0] in448;
input [7:0] in449;
input [7:0] in450;
input [7:0] in451;
input [7:0] in452;
input [7:0] in453;
input [7:0] in454;
input [7:0] in455;
input [7:0] in456;
input [7:0] in457;
input [7:0] in458;
input [7:0] in459;
input [7:0] in460;
input [7:0] in461;
input [7:0] in462;
input [7:0] in463;
input [7:0] in464;
input [7:0] in465;
input [7:0] in466;
input [7:0] in467;
input [7:0] in468;
input [7:0] in469;
input [7:0] in470;
input [7:0] in471;
input [7:0] in472;
input [7:0] in473;
input [7:0] in474;
input [7:0] in475;
input [7:0] in476;
input [7:0] in477;
input [7:0] in478;
input [7:0] in479;
input [7:0] in480;
input [7:0] in481;
input [7:0] in482;
input [7:0] in483;
input [7:0] in484;
input [7:0] in485;
input [7:0] in486;
input [7:0] in487;
input [7:0] in488;
input [7:0] in489;
input [7:0] in490;
input [7:0] in491;
input [7:0] in492;
input [7:0] in493;
input [7:0] in494;
input [7:0] in495;
input [7:0] in496;
input [7:0] in497;
input [7:0] in498;
input [7:0] in499;
input [7:0] in500;
input [7:0] in501;
input [7:0] in502;
input [7:0] in503;
input [7:0] in504;
input [7:0] in505;
input [7:0] in506;
input [7:0] in507;
input [7:0] in508;
input [7:0] in509;
input [7:0] in510;
input [7:0] in511;
input [7:0] in512;
input [7:0] in513;
input [7:0] in514;
input [7:0] in515;
input [7:0] in516;
input [7:0] in517;
input [7:0] in518;
input [7:0] in519;
input [7:0] in520;
input [7:0] in521;
input [7:0] in522;
input [7:0] in523;
input [7:0] in524;
input [7:0] in525;
input [7:0] in526;
input [7:0] in527;
input [7:0] in528;
input [7:0] in529;
input [7:0] in530;
input [7:0] in531;
input [7:0] in532;
input [7:0] in533;
input [7:0] in534;
input [7:0] in535;
input [7:0] in536;
input [7:0] in537;
input [7:0] in538;
input [7:0] in539;
input [7:0] in540;
input [7:0] in541;
input [7:0] in542;
input [7:0] in543;
input [7:0] in544;
input [7:0] in545;
input [7:0] in546;
input [7:0] in547;
input [7:0] in548;
input [7:0] in549;
input [7:0] in550;
input [7:0] in551;
input [7:0] in552;
input [7:0] in553;
input [7:0] in554;
input [7:0] in555;
input [7:0] in556;
input [7:0] in557;
input [7:0] in558;
input [7:0] in559;
input [7:0] in560;
input [7:0] in561;
input [7:0] in562;
input [7:0] in563;
input [7:0] in564;
input [7:0] in565;
input [7:0] in566;
input [7:0] in567;
input [7:0] in568;
input [7:0] in569;
input [7:0] in570;
input [7:0] in571;
input [7:0] in572;
input [7:0] in573;
input [7:0] in574;
input [7:0] in575;


 output [7:0] out0;
output [7:0] out1;
output [7:0] out2;
output [7:0] out3;
output [7:0] out4;
output [7:0] out5;
output [7:0] out6;
output [7:0] out7;
output [7:0] out8;
output [7:0] out9;
output [7:0] out10;
output [7:0] out11;
output [7:0] out12;
output [7:0] out13;
output [7:0] out14;
output [7:0] out15;
output [7:0] out16;
output [7:0] out17;
output [7:0] out18;
output [7:0] out19;
output [7:0] out20;
output [7:0] out21;
output [7:0] out22;
output [7:0] out23;
output [7:0] out24;
output [7:0] out25;
output [7:0] out26;
output [7:0] out27;
output [7:0] out28;
output [7:0] out29;
output [7:0] out30;
output [7:0] out31;
output [7:0] out32;
output [7:0] out33;
output [7:0] out34;
output [7:0] out35;
output [7:0] out36;
output [7:0] out37;
output [7:0] out38;
output [7:0] out39;
output [7:0] out40;
output [7:0] out41;
output [7:0] out42;
output [7:0] out43;
output [7:0] out44;
output [7:0] out45;
output [7:0] out46;
output [7:0] out47;
output [7:0] out48;
output [7:0] out49;
output [7:0] out50;
output [7:0] out51;
output [7:0] out52;
output [7:0] out53;
output [7:0] out54;
output [7:0] out55;
output [7:0] out56;
output [7:0] out57;
output [7:0] out58;
output [7:0] out59;
output [7:0] out60;
output [7:0] out61;
output [7:0] out62;
output [7:0] out63;
output [7:0] out64;
output [7:0] out65;
output [7:0] out66;
output [7:0] out67;
output [7:0] out68;
output [7:0] out69;
output [7:0] out70;
output [7:0] out71;
output [7:0] out72;
output [7:0] out73;
output [7:0] out74;
output [7:0] out75;
output [7:0] out76;
output [7:0] out77;
output [7:0] out78;
output [7:0] out79;
output [7:0] out80;
output [7:0] out81;
output [7:0] out82;
output [7:0] out83;
output [7:0] out84;
output [7:0] out85;
output [7:0] out86;
output [7:0] out87;
output [7:0] out88;
output [7:0] out89;
output [7:0] out90;
output [7:0] out91;
output [7:0] out92;
output [7:0] out93;
output [7:0] out94;
output [7:0] out95;
output [7:0] out96;
output [7:0] out97;
output [7:0] out98;
output [7:0] out99;
output [7:0] out100;
output [7:0] out101;
output [7:0] out102;
output [7:0] out103;
output [7:0] out104;
output [7:0] out105;
output [7:0] out106;
output [7:0] out107;
output [7:0] out108;
output [7:0] out109;
output [7:0] out110;
output [7:0] out111;
output [7:0] out112;
output [7:0] out113;
output [7:0] out114;
output [7:0] out115;
output [7:0] out116;
output [7:0] out117;
output [7:0] out118;
output [7:0] out119;
output [7:0] out120;
output [7:0] out121;
output [7:0] out122;
output [7:0] out123;
output [7:0] out124;
output [7:0] out125;
output [7:0] out126;
output [7:0] out127;
output [7:0] out128;
output [7:0] out129;
output [7:0] out130;
output [7:0] out131;
output [7:0] out132;
output [7:0] out133;
output [7:0] out134;
output [7:0] out135;
output [7:0] out136;
output [7:0] out137;
output [7:0] out138;
output [7:0] out139;
output [7:0] out140;
output [7:0] out141;
output [7:0] out142;
output [7:0] out143;
output ready;


pooling_dp dp1( .in0(in0),.in1(in1),.in2(in2),.in3(in3),.in4(in4),.in5(in5),.in6(in6),.in7(in7),.in8(in8),.in9(in9),.in10(in10),.in11(in11),.in12(in12),.in13(in13),.in14(in14),.in15(in15),.in16(in16),.in17(in17),.in18(in18),.in19(in19),.in20(in20),.in21(in21),.in22(in22),.in23(in23),.in24(in24),.in25(in25),.in26(in26),.in27(in27),.in28(in28),.in29(in29),.in30(in30),.in31(in31),.in32(in32),.in33(in33),.in34(in34),.in35(in35),.in36(in36),.in37(in37),.in38(in38),.in39(in39),.in40(in40),.in41(in41),.in42(in42),.in43(in43),.in44(in44),.in45(in45),.in46(in46),.in47(in47),.in48(in48),.in49(in49),.in50(in50),.in51(in51),.in52(in52),.in53(in53),.in54(in54),.in55(in55),.in56(in56),.in57(in57),.in58(in58),.in59(in59),.in60(in60),.in61(in61),.in62(in62),.in63(in63),.in64(in64),.in65(in65),.in66(in66),.in67(in67),.in68(in68),.in69(in69),.in70(in70),.in71(in71),.in72(in72),.in73(in73),.in74(in74),.in75(in75),.in76(in76),.in77(in77),.in78(in78),.in79(in79),.in80(in80),.in81(in81),.in82(in82),.in83(in83),.in84(in84),.in85(in85),.in86(in86),.in87(in87),.in88(in88),.in89(in89),.in90(in90),.in91(in91),.in92(in92),.in93(in93),.in94(in94),.in95(in95),.in96(in96),.in97(in97),.in98(in98),.in99(in99),.in100(in100),.in101(in101),.in102(in102),.in103(in103),.in104(in104),.in105(in105),.in106(in106),.in107(in107),.in108(in108),.in109(in109),.in110(in110),.in111(in111),.in112(in112),.in113(in113),.in114(in114),.in115(in115),.in116(in116),.in117(in117),.in118(in118),.in119(in119),.in120(in120),.in121(in121),.in122(in122),.in123(in123),.in124(in124),.in125(in125),.in126(in126),.in127(in127),.in128(in128),.in129(in129),.in130(in130),.in131(in131),.in132(in132),.in133(in133),.in134(in134),.in135(in135),.in136(in136),.in137(in137),.in138(in138),.in139(in139),.in140(in140),.in141(in141),.in142(in142),.in143(in143),.in144(in144),.in145(in145),.in146(in146),.in147(in147),.in148(in148),.in149(in149),.in150(in150),.in151(in151),.in152(in152),.in153(in153),.in154(in154),.in155(in155),.in156(in156),.in157(in157),.in158(in158),.in159(in159),.in160(in160),.in161(in161),.in162(in162),.in163(in163),.in164(in164),.in165(in165),.in166(in166),.in167(in167),.in168(in168),.in169(in169),.in170(in170),.in171(in171),.in172(in172),.in173(in173),.in174(in174),.in175(in175),.in176(in176),.in177(in177),.in178(in178),.in179(in179),.in180(in180),.in181(in181),.in182(in182),.in183(in183),.in184(in184),.in185(in185),.in186(in186),.in187(in187),.in188(in188),.in189(in189),.in190(in190),.in191(in191),.in192(in192),.in193(in193),.in194(in194),.in195(in195),.in196(in196),.in197(in197),.in198(in198),.in199(in199),.in200(in200),.in201(in201),.in202(in202),.in203(in203),.in204(in204),.in205(in205),.in206(in206),.in207(in207),.in208(in208),.in209(in209),.in210(in210),.in211(in211),.in212(in212),.in213(in213),.in214(in214),.in215(in215),.in216(in216),.in217(in217),.in218(in218),.in219(in219),.in220(in220),.in221(in221),.in222(in222),.in223(in223),.in224(in224),.in225(in225),.in226(in226),.in227(in227),.in228(in228),.in229(in229),.in230(in230),.in231(in231),.in232(in232),.in233(in233),.in234(in234),.in235(in235),.in236(in236),.in237(in237),.in238(in238),.in239(in239),.in240(in240),.in241(in241),.in242(in242),.in243(in243),.in244(in244),.in245(in245),.in246(in246),.in247(in247),.in248(in248),.in249(in249),.in250(in250),.in251(in251),.in252(in252),.in253(in253),.in254(in254),.in255(in255),.in256(in256),.in257(in257),.in258(in258),.in259(in259),.in260(in260),.in261(in261),.in262(in262),.in263(in263),.in264(in264),.in265(in265),.in266(in266),.in267(in267),.in268(in268),.in269(in269),.in270(in270),.in271(in271),.in272(in272),.in273(in273),.in274(in274),.in275(in275),.in276(in276),.in277(in277),.in278(in278),.in279(in279),.in280(in280),.in281(in281),.in282(in282),.in283(in283),.in284(in284),.in285(in285),.in286(in286),.in287(in287),.in288(in288),.in289(in289),.in290(in290),.in291(in291),.in292(in292),.in293(in293),.in294(in294),.in295(in295),.in296(in296),.in297(in297),.in298(in298),.in299(in299),.in300(in300),.in301(in301),.in302(in302),.in303(in303),.in304(in304),.in305(in305),.in306(in306),.in307(in307),.in308(in308),.in309(in309),.in310(in310),.in311(in311),.in312(in312),.in313(in313),.in314(in314),.in315(in315),.in316(in316),.in317(in317),.in318(in318),.in319(in319),.in320(in320),.in321(in321),.in322(in322),.in323(in323),.in324(in324),.in325(in325),.in326(in326),.in327(in327),.in328(in328),.in329(in329),.in330(in330),.in331(in331),.in332(in332),.in333(in333),.in334(in334),.in335(in335),.in336(in336),.in337(in337),.in338(in338),.in339(in339),.in340(in340),.in341(in341),.in342(in342),.in343(in343),.in344(in344),.in345(in345),.in346(in346),.in347(in347),.in348(in348),.in349(in349),.in350(in350),.in351(in351),.in352(in352),.in353(in353),.in354(in354),.in355(in355),.in356(in356),.in357(in357),.in358(in358),.in359(in359),.in360(in360),.in361(in361),.in362(in362),.in363(in363),.in364(in364),.in365(in365),.in366(in366),.in367(in367),.in368(in368),.in369(in369),.in370(in370),.in371(in371),.in372(in372),.in373(in373),.in374(in374),.in375(in375),.in376(in376),.in377(in377),.in378(in378),.in379(in379),.in380(in380),.in381(in381),.in382(in382),.in383(in383),.in384(in384),.in385(in385),.in386(in386),.in387(in387),.in388(in388),.in389(in389),.in390(in390),.in391(in391),.in392(in392),.in393(in393),.in394(in394),.in395(in395),.in396(in396),.in397(in397),.in398(in398),.in399(in399),.in400(in400),.in401(in401),.in402(in402),.in403(in403),.in404(in404),.in405(in405),.in406(in406),.in407(in407),.in408(in408),.in409(in409),.in410(in410),.in411(in411),.in412(in412),.in413(in413),.in414(in414),.in415(in415),.in416(in416),.in417(in417),.in418(in418),.in419(in419),.in420(in420),.in421(in421),.in422(in422),.in423(in423),.in424(in424),.in425(in425),.in426(in426),.in427(in427),.in428(in428),.in429(in429),.in430(in430),.in431(in431),.in432(in432),.in433(in433),.in434(in434),.in435(in435),.in436(in436),.in437(in437),.in438(in438),.in439(in439),.in440(in440),.in441(in441),.in442(in442),.in443(in443),.in444(in444),.in445(in445),.in446(in446),.in447(in447),.in448(in448),.in449(in449),.in450(in450),.in451(in451),.in452(in452),.in453(in453),.in454(in454),.in455(in455),.in456(in456),.in457(in457),.in458(in458),.in459(in459),.in460(in460),.in461(in461),.in462(in462),.in463(in463),.in464(in464),.in465(in465),.in466(in466),.in467(in467),.in468(in468),.in469(in469),.in470(in470),.in471(in471),.in472(in472),.in473(in473),.in474(in474),.in475(in475),.in476(in476),.in477(in477),.in478(in478),.in479(in479),.in480(in480),.in481(in481),.in482(in482),.in483(in483),.in484(in484),.in485(in485),.in486(in486),.in487(in487),.in488(in488),.in489(in489),.in490(in490),.in491(in491),.in492(in492),.in493(in493),.in494(in494),.in495(in495),.in496(in496),.in497(in497),.in498(in498),.in499(in499),.in500(in500),.in501(in501),.in502(in502),.in503(in503),.in504(in504),.in505(in505),.in506(in506),.in507(in507),.in508(in508),.in509(in509),.in510(in510),.in511(in511),.in512(in512),.in513(in513),.in514(in514),.in515(in515),.in516(in516),.in517(in517),.in518(in518),.in519(in519),.in520(in520),.in521(in521),.in522(in522),.in523(in523),.in524(in524),.in525(in525),.in526(in526),.in527(in527),.in528(in528),.in529(in529),.in530(in530),.in531(in531),.in532(in532),.in533(in533),.in534(in534),.in535(in535),.in536(in536),.in537(in537),.in538(in538),.in539(in539),.in540(in540),.in541(in541),.in542(in542),.in543(in543),.in544(in544),.in545(in545),.in546(in546),.in547(in547),.in548(in548),.in549(in549),.in550(in550),.in551(in551),.in552(in552),.in553(in553),.in554(in554),.in555(in555),.in556(in556),.in557(in557),.in558(in558),.in559(in559),.in560(in560),.in561(in561),.in562(in562),.in563(in563),.in564(in564),.in565(in565),.in566(in566),.in567(in567),.in568(in568),.in569(in569),.in570(in570),.in571(in571),.in572(in572),.in573(in573),.in574(in574),.in575(in575),
 .out0(out0),.out1(out1),.out2(out2),.out3(out3),.out4(out4),.out5(out5),.out6(out6),.out7(out7),.out8(out8),.out9(out9),.out10(out10),.out11(out11),.out12(out12),.out13(out13),.out14(out14),.out15(out15),.out16(out16),.out17(out17),.out18(out18),.out19(out19),.out20(out20),.out21(out21),.out22(out22),.out23(out23),.out24(out24),.out25(out25),.out26(out26),.out27(out27),.out28(out28),.out29(out29),.out30(out30),.out31(out31),.out32(out32),.out33(out33),.out34(out34),.out35(out35),.out36(out36),.out37(out37),.out38(out38),.out39(out39),.out40(out40),.out41(out41),.out42(out42),.out43(out43),.out44(out44),.out45(out45),.out46(out46),.out47(out47),.out48(out48),.out49(out49),.out50(out50),.out51(out51),.out52(out52),.out53(out53),.out54(out54),.out55(out55),.out56(out56),.out57(out57),.out58(out58),.out59(out59),.out60(out60),.out61(out61),.out62(out62),.out63(out63),.out64(out64),.out65(out65),.out66(out66),.out67(out67),.out68(out68),.out69(out69),.out70(out70),.out71(out71),.out72(out72),.out73(out73),.out74(out74),.out75(out75),.out76(out76),.out77(out77),.out78(out78),.out79(out79),.out80(out80),.out81(out81),.out82(out82),.out83(out83),.out84(out84),.out85(out85),.out86(out86),.out87(out87),.out88(out88),.out89(out89),.out90(out90),.out91(out91),.out92(out92),.out93(out93),.out94(out94),.out95(out95),.out96(out96),.out97(out97),.out98(out98),.out99(out99),.out100(out100),.out101(out101),.out102(out102),.out103(out103),.out104(out104),.out105(out105),.out106(out106),.out107(out107),.out108(out108),.out109(out109),.out110(out110),.out111(out111),.out112(out112),.out113(out113),.out114(out114),.out115(out115),.out116(out116),.out117(out117),.out118(out118),.out119(out119),.out120(out120),.out121(out121),.out122(out122),.out123(out123),.out124(out124),.out125(out125),.out126(out126),.out127(out127),.out128(out128),.out129(out129),.out130(out130),.out131(out131),.out132(out132),.out133(out133),.out134(out134),.out135(out135),.out136(out136),.out137(out137),.out138(out138),.out139(out139),.out140(out140),.out141(out141),.out142(out142),.out143(out143)
 ,.ready(ready),.clk(clk),.start(start));
 


endmodule



module pooling_dp(in0,in1,in2,in3,in4,in5,in6,in7,in8,in9,in10,in11,in12,in13,in14,
in15,in16,in17,in18,in19,in20,in21,in22,in23,in24,in25,in26,in27,in28,in29,in30,in31,
in32,in33,in34,in35,in36,in37,in38,in39,in40,in41,in42,in43,in44,in45,in46,in47,in48,
in49,in50,in51,in52,in53,in54,in55,in56,in57,in58,in59,in60,in61,in62,in63,in64,in65,
in66,in67,in68,in69,in70,in71,in72,in73,in74,in75,in76,in77,in78,in79,in80,in81,in82,
in83,in84,in85,in86,in87,in88,in89,in90,in91,in92,in93,in94,in95,in96,in97,in98,in99,
in100,in101,in102,in103,in104,in105,in106,in107,in108,in109,in110,in111,in112,in113,
in114,in115,in116,in117,in118,in119,in120,in121,in122,in123,in124,in125,in126,in127,
in128,in129,in130,in131,in132,in133,in134,in135,in136,in137,in138,in139,in140,in141,
in142,in143,in144,in145,in146,in147,in148,in149,in150,in151,in152,in153,in154,in155,
in156,in157,in158,in159,in160,in161,in162,in163,in164,in165,in166,in167,in168,in169,
in170,in171,in172,in173,in174,in175,in176,in177,in178,in179,in180,in181,in182,in183,
in184,in185,in186,in187,in188,in189,in190,in191,in192,in193,in194,in195,in196,in197,
in198,in199,in200,in201,in202,in203,in204,in205,in206,in207,in208,in209,in210,in211,
in212,in213,in214,in215,in216,in217,in218,in219,in220,in221,in222,in223,in224,in225,
in226,in227,in228,in229,in230,in231,in232,in233,in234,in235,in236,in237,in238,in239,
in240,in241,in242,in243,in244,in245,in246,in247,in248,in249,in250,in251,in252,in253,
in254,in255,in256,in257,in258,in259,in260,in261,in262,in263,in264,in265,in266,in267,
in268,in269,in270,in271,in272,in273,in274,in275,in276,in277,in278,in279,in280,in281,
in282,in283,in284,in285,in286,in287,in288,in289,in290,in291,in292,in293,in294,in295,
in296,in297,in298,in299,in300,in301,in302,in303,in304,in305,in306,in307,in308,in309,
in310,in311,in312,in313,in314,in315,in316,in317,in318,in319,in320,in321,in322,in323,
in324,in325,in326,in327,in328,in329,in330,in331,in332,in333,in334,in335,in336,in337,
in338,in339,in340,in341,in342,in343,in344,in345,in346,in347,in348,in349,in350,in351,
in352,in353,in354,in355,in356,in357,in358,in359,in360,in361,in362,in363,in364,in365,in366,
in367,in368,in369,in370,in371,in372,in373,in374,in375,in376,in377,in378,in379,in380,
in381,in382,in383,in384,in385,in386,in387,in388,in389,in390,in391,in392,in393,in394,
in395,in396,in397,in398,in399,in400,in401,in402,in403,in404,in405,in406,in407,in408,
in409,in410,in411,in412,in413,in414,in415,in416,in417,in418,in419,in420,in421,in422,
in423,in424,in425,in426,in427,in428,in429,in430,in431,in432,in433,in434,in435,in436,
in437,in438,in439,in440,in441,in442,in443,in444,in445,in446,in447,in448,in449,in450,
in451,in452,in453,in454,in455,in456,in457,in458,in459,in460,in461,in462,in463,in464,
in465,in466,in467,in468,in469,in470,in471,in472,in473,in474,in475,in476,in477,in478,
in479,in480,in481,in482,in483,in484,in485,in486,in487,in488,in489,in490,in491,in492,
in493,in494,in495,in496,in497,in498,in499,in500,in501,in502,in503,in504,in505,in506,
in507,in508,in509,in510,in511,in512,in513,in514,in515,in516,in517,in518,in519,in520,
in521,in522,in523,in524,in525,in526,in527,in528,in529,in530,in531,in532,in533,in534,
in535,in536,in537,in538,in539,in540,in541,in542,in543,in544,in545,in546,in547,in548,
in549,in550,in551,in552,in553,in554,in555,in556,in557,in558,in559,in560,in561,in562,
in563,in564,in565,in566,in567,in568,in569,in570,in571,in572,in573,in574,in575,out0,out1,out2,out3,out4,out5,out6,out7,out8,out9,out10,out11,out12,out13,out14,out15,out16,out17,out18,out19,out20,out21,out22,out23,out24,out25,out26,out27,out28,out29,out30,out31,out32,out33,out34,out35,out36,out37,out38,out39,out40,out41,out42,out43,out44,out45,out46,out47,out48,out49,out50,out51,out52,out53,out54,out55,out56,out57,out58,out59,out60,out61,out62,out63,out64,out65,out66,out67,out68,out69,out70,out71,out72,out73,out74,out75,out76,out77,out78,out79,out80,out81,out82,out83,out84,out85,out86,out87,out88,out89,out90,out91,out92,out93,out94,out95,out96,out97,out98,out99,out100,out101,out102,out103,out104,out105,out106,out107,out108,out109,out110,out111,out112,out113,out114,out115,out116,out117,out118,out119,out120,out121,out122,out123,out124,out125,out126,out127,out128,out129,out130,out131,out132,out133,out134,out135,out136,out137,out138,out139,out140,out141,out142,out143,
clk,start,ready);

input clk;
input start;
input [7:0] in0;
input [7:0] in1;
input [7:0] in2;
input [7:0] in3;
input [7:0] in4;
input [7:0] in5;
input [7:0] in6;
input [7:0] in7;
input [7:0] in8;
input [7:0] in9;
input [7:0] in10;
input [7:0] in11;
input [7:0] in12;
input [7:0] in13;
input [7:0] in14;
input [7:0] in15;
input [7:0] in16;
input [7:0] in17;
input [7:0] in18;
input [7:0] in19;
input [7:0] in20;
input [7:0] in21;
input [7:0] in22;
input [7:0] in23;
input [7:0] in24;
input [7:0] in25;
input [7:0] in26;
input [7:0] in27;
input [7:0] in28;
input [7:0] in29;
input [7:0] in30;
input [7:0] in31;
input [7:0] in32;
input [7:0] in33;
input [7:0] in34;
input [7:0] in35;
input [7:0] in36;
input [7:0] in37;
input [7:0] in38;
input [7:0] in39;
input [7:0] in40;
input [7:0] in41;
input [7:0] in42;
input [7:0] in43;
input [7:0] in44;
input [7:0] in45;
input [7:0] in46;
input [7:0] in47;
input [7:0] in48;
input [7:0] in49;
input [7:0] in50;
input [7:0] in51;
input [7:0] in52;
input [7:0] in53;
input [7:0] in54;
input [7:0] in55;
input [7:0] in56;
input [7:0] in57;
input [7:0] in58;
input [7:0] in59;
input [7:0] in60;
input [7:0] in61;
input [7:0] in62;
input [7:0] in63;
input [7:0] in64;
input [7:0] in65;
input [7:0] in66;
input [7:0] in67;
input [7:0] in68;
input [7:0] in69;
input [7:0] in70;
input [7:0] in71;
input [7:0] in72;
input [7:0] in73;
input [7:0] in74;
input [7:0] in75;
input [7:0] in76;
input [7:0] in77;
input [7:0] in78;
input [7:0] in79;
input [7:0] in80;
input [7:0] in81;
input [7:0] in82;
input [7:0] in83;
input [7:0] in84;
input [7:0] in85;
input [7:0] in86;
input [7:0] in87;
input [7:0] in88;
input [7:0] in89;
input [7:0] in90;
input [7:0] in91;
input [7:0] in92;
input [7:0] in93;
input [7:0] in94;
input [7:0] in95;
input [7:0] in96;
input [7:0] in97;
input [7:0] in98;
input [7:0] in99;
input [7:0] in100;
input [7:0] in101;
input [7:0] in102;
input [7:0] in103;
input [7:0] in104;
input [7:0] in105;
input [7:0] in106;
input [7:0] in107;
input [7:0] in108;
input [7:0] in109;
input [7:0] in110;
input [7:0] in111;
input [7:0] in112;
input [7:0] in113;
input [7:0] in114;
input [7:0] in115;
input [7:0] in116;
input [7:0] in117;
input [7:0] in118;
input [7:0] in119;
input [7:0] in120;
input [7:0] in121;
input [7:0] in122;
input [7:0] in123;
input [7:0] in124;
input [7:0] in125;
input [7:0] in126;
input [7:0] in127;
input [7:0] in128;
input [7:0] in129;
input [7:0] in130;
input [7:0] in131;
input [7:0] in132;
input [7:0] in133;
input [7:0] in134;
input [7:0] in135;
input [7:0] in136;
input [7:0] in137;
input [7:0] in138;
input [7:0] in139;
input [7:0] in140;
input [7:0] in141;
input [7:0] in142;
input [7:0] in143;
input [7:0] in144;
input [7:0] in145;
input [7:0] in146;
input [7:0] in147;
input [7:0] in148;
input [7:0] in149;
input [7:0] in150;
input [7:0] in151;
input [7:0] in152;
input [7:0] in153;
input [7:0] in154;
input [7:0] in155;
input [7:0] in156;
input [7:0] in157;
input [7:0] in158;
input [7:0] in159;
input [7:0] in160;
input [7:0] in161;
input [7:0] in162;
input [7:0] in163;
input [7:0] in164;
input [7:0] in165;
input [7:0] in166;
input [7:0] in167;
input [7:0] in168;
input [7:0] in169;
input [7:0] in170;
input [7:0] in171;
input [7:0] in172;
input [7:0] in173;
input [7:0] in174;
input [7:0] in175;
input [7:0] in176;
input [7:0] in177;
input [7:0] in178;
input [7:0] in179;
input [7:0] in180;
input [7:0] in181;
input [7:0] in182;
input [7:0] in183;
input [7:0] in184;
input [7:0] in185;
input [7:0] in186;
input [7:0] in187;
input [7:0] in188;
input [7:0] in189;
input [7:0] in190;
input [7:0] in191;
input [7:0] in192;
input [7:0] in193;
input [7:0] in194;
input [7:0] in195;
input [7:0] in196;
input [7:0] in197;
input [7:0] in198;
input [7:0] in199;
input [7:0] in200;
input [7:0] in201;
input [7:0] in202;
input [7:0] in203;
input [7:0] in204;
input [7:0] in205;
input [7:0] in206;
input [7:0] in207;
input [7:0] in208;
input [7:0] in209;
input [7:0] in210;
input [7:0] in211;
input [7:0] in212;
input [7:0] in213;
input [7:0] in214;
input [7:0] in215;
input [7:0] in216;
input [7:0] in217;
input [7:0] in218;
input [7:0] in219;
input [7:0] in220;
input [7:0] in221;
input [7:0] in222;
input [7:0] in223;
input [7:0] in224;
input [7:0] in225;
input [7:0] in226;
input [7:0] in227;
input [7:0] in228;
input [7:0] in229;
input [7:0] in230;
input [7:0] in231;
input [7:0] in232;
input [7:0] in233;
input [7:0] in234;
input [7:0] in235;
input [7:0] in236;
input [7:0] in237;
input [7:0] in238;
input [7:0] in239;
input [7:0] in240;
input [7:0] in241;
input [7:0] in242;
input [7:0] in243;
input [7:0] in244;
input [7:0] in245;
input [7:0] in246;
input [7:0] in247;
input [7:0] in248;
input [7:0] in249;
input [7:0] in250;
input [7:0] in251;
input [7:0] in252;
input [7:0] in253;
input [7:0] in254;
input [7:0] in255;
input [7:0] in256;
input [7:0] in257;
input [7:0] in258;
input [7:0] in259;
input [7:0] in260;
input [7:0] in261;
input [7:0] in262;
input [7:0] in263;
input [7:0] in264;
input [7:0] in265;
input [7:0] in266;
input [7:0] in267;
input [7:0] in268;
input [7:0] in269;
input [7:0] in270;
input [7:0] in271;
input [7:0] in272;
input [7:0] in273;
input [7:0] in274;
input [7:0] in275;
input [7:0] in276;
input [7:0] in277;
input [7:0] in278;
input [7:0] in279;
input [7:0] in280;
input [7:0] in281;
input [7:0] in282;
input [7:0] in283;
input [7:0] in284;
input [7:0] in285;
input [7:0] in286;
input [7:0] in287;
input [7:0] in288;
input [7:0] in289;
input [7:0] in290;
input [7:0] in291;
input [7:0] in292;
input [7:0] in293;
input [7:0] in294;
input [7:0] in295;
input [7:0] in296;
input [7:0] in297;
input [7:0] in298;
input [7:0] in299;
input [7:0] in300;
input [7:0] in301;
input [7:0] in302;
input [7:0] in303;
input [7:0] in304;
input [7:0] in305;
input [7:0] in306;
input [7:0] in307;
input [7:0] in308;
input [7:0] in309;
input [7:0] in310;
input [7:0] in311;
input [7:0] in312;
input [7:0] in313;
input [7:0] in314;
input [7:0] in315;
input [7:0] in316;
input [7:0] in317;
input [7:0] in318;
input [7:0] in319;
input [7:0] in320;
input [7:0] in321;
input [7:0] in322;
input [7:0] in323;
input [7:0] in324;
input [7:0] in325;
input [7:0] in326;
input [7:0] in327;
input [7:0] in328;
input [7:0] in329;
input [7:0] in330;
input [7:0] in331;
input [7:0] in332;
input [7:0] in333;
input [7:0] in334;
input [7:0] in335;
input [7:0] in336;
input [7:0] in337;
input [7:0] in338;
input [7:0] in339;
input [7:0] in340;
input [7:0] in341;
input [7:0] in342;
input [7:0] in343;
input [7:0] in344;
input [7:0] in345;
input [7:0] in346;
input [7:0] in347;
input [7:0] in348;
input [7:0] in349;
input [7:0] in350;
input [7:0] in351;
input [7:0] in352;
input [7:0] in353;
input [7:0] in354;
input [7:0] in355;
input [7:0] in356;
input [7:0] in357;
input [7:0] in358;
input [7:0] in359;
input [7:0] in360;
input [7:0] in361;
input [7:0] in362;
input [7:0] in363;
input [7:0] in364;
input [7:0] in365;
input [7:0] in366;
input [7:0] in367;
input [7:0] in368;
input [7:0] in369;
input [7:0] in370;
input [7:0] in371;
input [7:0] in372;
input [7:0] in373;
input [7:0] in374;
input [7:0] in375;
input [7:0] in376;
input [7:0] in377;
input [7:0] in378;
input [7:0] in379;
input [7:0] in380;
input [7:0] in381;
input [7:0] in382;
input [7:0] in383;
input [7:0] in384;
input [7:0] in385;
input [7:0] in386;
input [7:0] in387;
input [7:0] in388;
input [7:0] in389;
input [7:0] in390;
input [7:0] in391;
input [7:0] in392;
input [7:0] in393;
input [7:0] in394;
input [7:0] in395;
input [7:0] in396;
input [7:0] in397;
input [7:0] in398;
input [7:0] in399;
input [7:0] in400;
input [7:0] in401;
input [7:0] in402;
input [7:0] in403;
input [7:0] in404;
input [7:0] in405;
input [7:0] in406;
input [7:0] in407;
input [7:0] in408;
input [7:0] in409;
input [7:0] in410;
input [7:0] in411;
input [7:0] in412;
input [7:0] in413;
input [7:0] in414;
input [7:0] in415;
input [7:0] in416;
input [7:0] in417;
input [7:0] in418;
input [7:0] in419;
input [7:0] in420;
input [7:0] in421;
input [7:0] in422;
input [7:0] in423;
input [7:0] in424;
input [7:0] in425;
input [7:0] in426;
input [7:0] in427;
input [7:0] in428;
input [7:0] in429;
input [7:0] in430;
input [7:0] in431;
input [7:0] in432;
input [7:0] in433;
input [7:0] in434;
input [7:0] in435;
input [7:0] in436;
input [7:0] in437;
input [7:0] in438;
input [7:0] in439;
input [7:0] in440;
input [7:0] in441;
input [7:0] in442;
input [7:0] in443;
input [7:0] in444;
input [7:0] in445;
input [7:0] in446;
input [7:0] in447;
input [7:0] in448;
input [7:0] in449;
input [7:0] in450;
input [7:0] in451;
input [7:0] in452;
input [7:0] in453;
input [7:0] in454;
input [7:0] in455;
input [7:0] in456;
input [7:0] in457;
input [7:0] in458;
input [7:0] in459;
input [7:0] in460;
input [7:0] in461;
input [7:0] in462;
input [7:0] in463;
input [7:0] in464;
input [7:0] in465;
input [7:0] in466;
input [7:0] in467;
input [7:0] in468;
input [7:0] in469;
input [7:0] in470;
input [7:0] in471;
input [7:0] in472;
input [7:0] in473;
input [7:0] in474;
input [7:0] in475;
input [7:0] in476;
input [7:0] in477;
input [7:0] in478;
input [7:0] in479;
input [7:0] in480;
input [7:0] in481;
input [7:0] in482;
input [7:0] in483;
input [7:0] in484;
input [7:0] in485;
input [7:0] in486;
input [7:0] in487;
input [7:0] in488;
input [7:0] in489;
input [7:0] in490;
input [7:0] in491;
input [7:0] in492;
input [7:0] in493;
input [7:0] in494;
input [7:0] in495;
input [7:0] in496;
input [7:0] in497;
input [7:0] in498;
input [7:0] in499;
input [7:0] in500;
input [7:0] in501;
input [7:0] in502;
input [7:0] in503;
input [7:0] in504;
input [7:0] in505;
input [7:0] in506;
input [7:0] in507;
input [7:0] in508;
input [7:0] in509;
input [7:0] in510;
input [7:0] in511;
input [7:0] in512;
input [7:0] in513;
input [7:0] in514;
input [7:0] in515;
input [7:0] in516;
input [7:0] in517;
input [7:0] in518;
input [7:0] in519;
input [7:0] in520;
input [7:0] in521;
input [7:0] in522;
input [7:0] in523;
input [7:0] in524;
input [7:0] in525;
input [7:0] in526;
input [7:0] in527;
input [7:0] in528;
input [7:0] in529;
input [7:0] in530;
input [7:0] in531;
input [7:0] in532;
input [7:0] in533;
input [7:0] in534;
input [7:0] in535;
input [7:0] in536;
input [7:0] in537;
input [7:0] in538;
input [7:0] in539;
input [7:0] in540;
input [7:0] in541;
input [7:0] in542;
input [7:0] in543;
input [7:0] in544;
input [7:0] in545;
input [7:0] in546;
input [7:0] in547;
input [7:0] in548;
input [7:0] in549;
input [7:0] in550;
input [7:0] in551;
input [7:0] in552;
input [7:0] in553;
input [7:0] in554;
input [7:0] in555;
input [7:0] in556;
input [7:0] in557;
input [7:0] in558;
input [7:0] in559;
input [7:0] in560;
input [7:0] in561;
input [7:0] in562;
input [7:0] in563;
input [7:0] in564;
input [7:0] in565;
input [7:0] in566;
input [7:0] in567;
input [7:0] in568;
input [7:0] in569;
input [7:0] in570;
input [7:0] in571;
input [7:0] in572;
input [7:0] in573;
input [7:0] in574;
input [7:0] in575;


 output [7:0] out0;
output [7:0] out1;
output [7:0] out2;
output [7:0] out3;
output [7:0] out4;
output [7:0] out5;
output [7:0] out6;
output [7:0] out7;
output [7:0] out8;
output [7:0] out9;
output [7:0] out10;
output [7:0] out11;
output [7:0] out12;
output [7:0] out13;
output [7:0] out14;
output [7:0] out15;
output [7:0] out16;
output [7:0] out17;
output [7:0] out18;
output [7:0] out19;
output [7:0] out20;
output [7:0] out21;
output [7:0] out22;
output [7:0] out23;
output [7:0] out24;
output [7:0] out25;
output [7:0] out26;
output [7:0] out27;
output [7:0] out28;
output [7:0] out29;
output [7:0] out30;
output [7:0] out31;
output [7:0] out32;
output [7:0] out33;
output [7:0] out34;
output [7:0] out35;
output [7:0] out36;
output [7:0] out37;
output [7:0] out38;
output [7:0] out39;
output [7:0] out40;
output [7:0] out41;
output [7:0] out42;
output [7:0] out43;
output [7:0] out44;
output [7:0] out45;
output [7:0] out46;
output [7:0] out47;
output [7:0] out48;
output [7:0] out49;
output [7:0] out50;
output [7:0] out51;
output [7:0] out52;
output [7:0] out53;
output [7:0] out54;
output [7:0] out55;
output [7:0] out56;
output [7:0] out57;
output [7:0] out58;
output [7:0] out59;
output [7:0] out60;
output [7:0] out61;
output [7:0] out62;
output [7:0] out63;
output [7:0] out64;
output [7:0] out65;
output [7:0] out66;
output [7:0] out67;
output [7:0] out68;
output [7:0] out69;
output [7:0] out70;
output [7:0] out71;
output [7:0] out72;
output [7:0] out73;
output [7:0] out74;
output [7:0] out75;
output [7:0] out76;
output [7:0] out77;
output [7:0] out78;
output [7:0] out79;
output [7:0] out80;
output [7:0] out81;
output [7:0] out82;
output [7:0] out83;
output [7:0] out84;
output [7:0] out85;
output [7:0] out86;
output [7:0] out87;
output [7:0] out88;
output [7:0] out89;
output [7:0] out90;
output [7:0] out91;
output [7:0] out92;
output [7:0] out93;
output [7:0] out94;
output [7:0] out95;
output [7:0] out96;
output [7:0] out97;
output [7:0] out98;
output [7:0] out99;
output [7:0] out100;
output [7:0] out101;
output [7:0] out102;
output [7:0] out103;
output [7:0] out104;
output [7:0] out105;
output [7:0] out106;
output [7:0] out107;
output [7:0] out108;
output [7:0] out109;
output [7:0] out110;
output [7:0] out111;
output [7:0] out112;
output [7:0] out113;
output [7:0] out114;
output [7:0] out115;
output [7:0] out116;
output [7:0] out117;
output [7:0] out118;
output [7:0] out119;
output [7:0] out120;
output [7:0] out121;
output [7:0] out122;
output [7:0] out123;
output [7:0] out124;
output [7:0] out125;
output [7:0] out126;
output [7:0] out127;
output [7:0] out128;
output [7:0] out129;
output [7:0] out130;
output [7:0] out131;
output [7:0] out132;
output [7:0] out133;
output [7:0] out134;
output [7:0] out135;
output [7:0] out136;
output [7:0] out137;
output [7:0] out138;
output [7:0] out139;
output [7:0] out140;
output [7:0] out141;
output [7:0] out142;
output [7:0] out143;
output ready;

 wire [7:0] muxpo0;
wire [7:0] muxpo1;
wire [7:0] muxpo2;
wire [7:0] muxpo3;
wire [7:0] muxpo4;
wire [7:0] muxpo5;
wire [7:0] muxpo6;
wire [7:0] muxpo7;
wire [7:0] muxpo8;
wire [7:0] muxpo9;
wire [7:0] muxpo10;
wire [7:0] muxpo11;
wire [7:0] muxpo12;
wire [7:0] muxpo13;
wire [7:0] muxpo14;
wire [7:0] muxpo15;
wire [7:0] muxpo16;
wire [7:0] muxpo17;
wire [7:0] muxpo18;
wire [7:0] muxpo19;
wire [7:0] muxpo20;
wire [7:0] muxpo21;
wire [7:0] muxpo22;
wire [7:0] muxpo23;
wire [7:0] muxpo24;
wire [7:0] muxpo25;
wire [7:0] muxpo26;
wire [7:0] muxpo27;
wire [7:0] muxpo28;
wire [7:0] muxpo29;
wire [7:0] muxpo30;
wire [7:0] muxpo31;
wire [7:0] muxpo32;
wire [7:0] muxpo33;
wire [7:0] muxpo34;
wire [7:0] muxpo35;
wire [7:0] muxpo36;
wire [7:0] muxpo37;
wire [7:0] muxpo38;
wire [7:0] muxpo39;
wire [7:0] muxpo40;
wire [7:0] muxpo41;
wire [7:0] muxpo42;
wire [7:0] muxpo43;
wire [7:0] muxpo44;
wire [7:0] muxpo45;
wire [7:0] muxpo46;
wire [7:0] muxpo47;
wire [7:0] muxpo48;
wire [7:0] muxpo49;
wire [7:0] muxpo50;
wire [7:0] muxpo51;
wire [7:0] muxpo52;
wire [7:0] muxpo53;
wire [7:0] muxpo54;
wire [7:0] muxpo55;
wire [7:0] muxpo56;
wire [7:0] muxpo57;
wire [7:0] muxpo58;
wire [7:0] muxpo59;
wire [7:0] muxpo60;
wire [7:0] muxpo61;
wire [7:0] muxpo62;
wire [7:0] muxpo63;
wire [7:0] muxpo64;
wire [7:0] muxpo65;
wire [7:0] muxpo66;
wire [7:0] muxpo67;
wire [7:0] muxpo68;
wire [7:0] muxpo69;
wire [7:0] muxpo70;
wire [7:0] muxpo71;
wire [7:0] muxpo72;
wire [7:0] muxpo73;
wire [7:0] muxpo74;
wire [7:0] muxpo75;
wire [7:0] muxpo76;
wire [7:0] muxpo77;
wire [7:0] muxpo78;
wire [7:0] muxpo79;
wire [7:0] muxpo80;
wire [7:0] muxpo81;
wire [7:0] muxpo82;
wire [7:0] muxpo83;
wire [7:0] muxpo84;
wire [7:0] muxpo85;
wire [7:0] muxpo86;
wire [7:0] muxpo87;
wire [7:0] muxpo88;
wire [7:0] muxpo89;
wire [7:0] muxpo90;
wire [7:0] muxpo91;
wire [7:0] muxpo92;
wire [7:0] muxpo93;
wire [7:0] muxpo94;
wire [7:0] muxpo95;
wire [7:0] muxpo96;
wire [7:0] muxpo97;
wire [7:0] muxpo98;
wire [7:0] muxpo99;
wire [7:0] muxpo100;
wire [7:0] muxpo101;
wire [7:0] muxpo102;
wire [7:0] muxpo103;
wire [7:0] muxpo104;
wire [7:0] muxpo105;
wire [7:0] muxpo106;
wire [7:0] muxpo107;
wire [7:0] muxpo108;
wire [7:0] muxpo109;
wire [7:0] muxpo110;
wire [7:0] muxpo111;
wire [7:0] muxpo112;
wire [7:0] muxpo113;
wire [7:0] muxpo114;
wire [7:0] muxpo115;
wire [7:0] muxpo116;
wire [7:0] muxpo117;
wire [7:0] muxpo118;
wire [7:0] muxpo119;
wire [7:0] muxpo120;
wire [7:0] muxpo121;
wire [7:0] muxpo122;
wire [7:0] muxpo123;
wire [7:0] muxpo124;
wire [7:0] muxpo125;
wire [7:0] muxpo126;
wire [7:0] muxpo127;
wire [7:0] muxpo128;
wire [7:0] muxpo129;
wire [7:0] muxpo130;
wire [7:0] muxpo131;
wire [7:0] muxpo132;
wire [7:0] muxpo133;
wire [7:0] muxpo134;
wire [7:0] muxpo135;
wire [7:0] muxpo136;
wire [7:0] muxpo137;
wire [7:0] muxpo138;
wire [7:0] muxpo139;
wire [7:0] muxpo140;
wire [7:0] muxpo141;
wire [7:0] muxpo142;
wire [7:0] muxpo143;

wire [7:0] muxpi0;wire [7:0] muxpi1;wire [7:0] muxpi2;wire [7:0] muxpi3;wire [7:0] muxpi4;wire [7:0] muxpi5;wire [7:0] muxpi6;wire [7:0] muxpi7;wire [7:0] muxpi8;wire [7:0] muxpi9;wire [7:0] muxpi10;wire [7:0] muxpi11;wire [7:0] muxpi12;wire [7:0] muxpi13;wire [7:0] muxpi14;wire [7:0] muxpi15;wire [7:0] muxpi16;wire [7:0] muxpi17;wire [7:0] muxpi18;wire [7:0] muxpi19;wire [7:0] muxpi20;wire [7:0] muxpi21;wire [7:0] muxpi22;wire [7:0] muxpi23;wire [7:0] muxpi24;wire [7:0] muxpi25;wire [7:0] muxpi26;wire [7:0] muxpi27;wire [7:0] muxpi28;wire [7:0] muxpi29;wire [7:0] muxpi30;wire [7:0] muxpi31;wire [7:0] muxpi32;wire [7:0] muxpi33;wire [7:0] muxpi34;wire [7:0] muxpi35;wire [7:0] muxpi36;wire [7:0] muxpi37;wire [7:0] muxpi38;wire [7:0] muxpi39;wire [7:0] muxpi40;wire [7:0] muxpi41;wire [7:0] muxpi42;wire [7:0] muxpi43;wire [7:0] muxpi44;wire [7:0] muxpi45;wire [7:0] muxpi46;wire [7:0] muxpi47;wire [7:0] muxpi48;wire [7:0] muxpi49;wire [7:0] muxpi50;wire [7:0] muxpi51;wire [7:0] muxpi52;wire [7:0] muxpi53;wire [7:0] muxpi54;wire [7:0] muxpi55;wire [7:0] muxpi56;wire [7:0] muxpi57;wire [7:0] muxpi58;wire [7:0] muxpi59;wire [7:0] muxpi60;wire [7:0] muxpi61;wire [7:0] muxpi62;wire [7:0] muxpi63;wire [7:0] muxpi64;wire [7:0] muxpi65;wire [7:0] muxpi66;wire [7:0] muxpi67;wire [7:0] muxpi68;wire [7:0] muxpi69;wire [7:0] muxpi70;wire [7:0] muxpi71;wire [7:0] muxpi72;wire [7:0] muxpi73;wire [7:0] muxpi74;wire [7:0] muxpi75;wire [7:0] muxpi76;wire [7:0] muxpi77;wire [7:0] muxpi78;wire [7:0] muxpi79;wire [7:0] muxpi80;wire [7:0] muxpi81;wire [7:0] muxpi82;wire [7:0] muxpi83;wire [7:0] muxpi84;wire [7:0] muxpi85;wire [7:0] muxpi86;wire [7:0] muxpi87;wire [7:0] muxpi88;wire [7:0] muxpi89;wire [7:0] muxpi90;wire [7:0] muxpi91;wire [7:0] muxpi92;wire [7:0] muxpi93;wire [7:0] muxpi94;wire [7:0] muxpi95;wire [7:0] muxpi96;wire [7:0] muxpi97;wire [7:0] muxpi98;wire [7:0] muxpi99;wire [7:0] muxpi100;wire [7:0] muxpi101;wire [7:0] muxpi102;wire [7:0] muxpi103;wire [7:0] muxpi104;wire [7:0] muxpi105;wire [7:0] muxpi106;wire [7:0] muxpi107;wire [7:0] muxpi108;wire [7:0] muxpi109;wire [7:0] muxpi110;wire [7:0] muxpi111;wire [7:0] muxpi112;wire [7:0] muxpi113;wire [7:0] muxpi114;wire [7:0] muxpi115;wire [7:0] muxpi116;wire [7:0] muxpi117;wire [7:0] muxpi118;wire [7:0] muxpi119;wire [7:0] muxpi120;wire [7:0] muxpi121;wire [7:0] muxpi122;wire [7:0] muxpi123;wire [7:0] muxpi124;wire [7:0] muxpi125;wire [7:0] muxpi126;wire [7:0] muxpi127;wire [7:0] muxpi128;wire [7:0] muxpi129;wire [7:0] muxpi130;wire [7:0] muxpi131;wire [7:0] muxpi132;wire [7:0] muxpi133;wire [7:0] muxpi134;wire [7:0] muxpi135;wire [7:0] muxpi136;wire [7:0] muxpi137;wire [7:0] muxpi138;wire [7:0] muxpi139;wire [7:0] muxpi140;wire [7:0] muxpi141;wire [7:0] muxpi142;wire [7:0] muxpi143;

 reg [7:0] muxreg0;
reg [7:0] muxreg1;
reg [7:0] muxreg2;
reg [7:0] muxreg3;
reg [7:0] muxreg4;
reg [7:0] muxreg5;
reg [7:0] muxreg6;
reg [7:0] muxreg7;
reg [7:0] muxreg8;
reg [7:0] muxreg9;
reg [7:0] muxreg10;
reg [7:0] muxreg11;
reg [7:0] muxreg12;
reg [7:0] muxreg13;
reg [7:0] muxreg14;
reg [7:0] muxreg15;
reg [7:0] muxreg16;
reg [7:0] muxreg17;
reg [7:0] muxreg18;
reg [7:0] muxreg19;
reg [7:0] muxreg20;
reg [7:0] muxreg21;
reg [7:0] muxreg22;
reg [7:0] muxreg23;
reg [7:0] muxreg24;
reg [7:0] muxreg25;
reg [7:0] muxreg26;
reg [7:0] muxreg27;
reg [7:0] muxreg28;
reg [7:0] muxreg29;
reg [7:0] muxreg30;
reg [7:0] muxreg31;
reg [7:0] muxreg32;
reg [7:0] muxreg33;
reg [7:0] muxreg34;
reg [7:0] muxreg35;
reg [7:0] muxreg36;
reg [7:0] muxreg37;
reg [7:0] muxreg38;
reg [7:0] muxreg39;
reg [7:0] muxreg40;
reg [7:0] muxreg41;
reg [7:0] muxreg42;
reg [7:0] muxreg43;
reg [7:0] muxreg44;
reg [7:0] muxreg45;
reg [7:0] muxreg46;
reg [7:0] muxreg47;
reg [7:0] muxreg48;
reg [7:0] muxreg49;
reg [7:0] muxreg50;
reg [7:0] muxreg51;
reg [7:0] muxreg52;
reg [7:0] muxreg53;
reg [7:0] muxreg54;
reg [7:0] muxreg55;
reg [7:0] muxreg56;
reg [7:0] muxreg57;
reg [7:0] muxreg58;
reg [7:0] muxreg59;
reg [7:0] muxreg60;
reg [7:0] muxreg61;
reg [7:0] muxreg62;
reg [7:0] muxreg63;
reg [7:0] muxreg64;
reg [7:0] muxreg65;
reg [7:0] muxreg66;
reg [7:0] muxreg67;
reg [7:0] muxreg68;
reg [7:0] muxreg69;
reg [7:0] muxreg70;
reg [7:0] muxreg71;
reg [7:0] muxreg72;
reg [7:0] muxreg73;
reg [7:0] muxreg74;
reg [7:0] muxreg75;
reg [7:0] muxreg76;
reg [7:0] muxreg77;
reg [7:0] muxreg78;
reg [7:0] muxreg79;
reg [7:0] muxreg80;
reg [7:0] muxreg81;
reg [7:0] muxreg82;
reg [7:0] muxreg83;
reg [7:0] muxreg84;
reg [7:0] muxreg85;
reg [7:0] muxreg86;
reg [7:0] muxreg87;
reg [7:0] muxreg88;
reg [7:0] muxreg89;
reg [7:0] muxreg90;
reg [7:0] muxreg91;
reg [7:0] muxreg92;
reg [7:0] muxreg93;
reg [7:0] muxreg94;
reg [7:0] muxreg95;
reg [7:0] muxreg96;
reg [7:0] muxreg97;
reg [7:0] muxreg98;
reg [7:0] muxreg99;
reg [7:0] muxreg100;
reg [7:0] muxreg101;
reg [7:0] muxreg102;
reg [7:0] muxreg103;
reg [7:0] muxreg104;
reg [7:0] muxreg105;
reg [7:0] muxreg106;
reg [7:0] muxreg107;
reg [7:0] muxreg108;
reg [7:0] muxreg109;
reg [7:0] muxreg110;
reg [7:0] muxreg111;
reg [7:0] muxreg112;
reg [7:0] muxreg113;
reg [7:0] muxreg114;
reg [7:0] muxreg115;
reg [7:0] muxreg116;
reg [7:0] muxreg117;
reg [7:0] muxreg118;
reg [7:0] muxreg119;
reg [7:0] muxreg120;
reg [7:0] muxreg121;
reg [7:0] muxreg122;
reg [7:0] muxreg123;
reg [7:0] muxreg124;
reg [7:0] muxreg125;
reg [7:0] muxreg126;
reg [7:0] muxreg127;
reg [7:0] muxreg128;
reg [7:0] muxreg129;
reg [7:0] muxreg130;
reg [7:0] muxreg131;
reg [7:0] muxreg132;
reg [7:0] muxreg133;
reg [7:0] muxreg134;
reg [7:0] muxreg135;
reg [7:0] muxreg136;
reg [7:0] muxreg137;
reg [7:0] muxreg138;
reg [7:0] muxreg139;
reg [7:0] muxreg140;
reg [7:0] muxreg141;
reg [7:0] muxreg142;
reg [7:0] muxreg143;

mux42 mux42p0(.a(in0),.b(in144),.c(in288),.d(in432),.sel(cs[1:0]),.out(muxpo0));
mux42 mux42p1(.a(in1),.b(in145),.c(in289),.d(in433),.sel(cs[1:0]),.out(muxpo1));
mux42 mux42p2(.a(in2),.b(in146),.c(in290),.d(in434),.sel(cs[1:0]),.out(muxpo2));
mux42 mux42p3(.a(in3),.b(in147),.c(in291),.d(in435),.sel(cs[1:0]),.out(muxpo3));
mux42 mux42p4(.a(in4),.b(in148),.c(in292),.d(in436),.sel(cs[1:0]),.out(muxpo4));
mux42 mux42p5(.a(in5),.b(in149),.c(in293),.d(in437),.sel(cs[1:0]),.out(muxpo5));
mux42 mux42p6(.a(in6),.b(in150),.c(in294),.d(in438),.sel(cs[1:0]),.out(muxpo6));
mux42 mux42p7(.a(in7),.b(in151),.c(in295),.d(in439),.sel(cs[1:0]),.out(muxpo7));
mux42 mux42p8(.a(in8),.b(in152),.c(in296),.d(in440),.sel(cs[1:0]),.out(muxpo8));
mux42 mux42p9(.a(in9),.b(in153),.c(in297),.d(in441),.sel(cs[1:0]),.out(muxpo9));
mux42 mux42p10(.a(in10),.b(in154),.c(in298),.d(in442),.sel(cs[1:0]),.out(muxpo10));
mux42 mux42p11(.a(in11),.b(in155),.c(in299),.d(in443),.sel(cs[1:0]),.out(muxpo11));
mux42 mux42p12(.a(in12),.b(in156),.c(in300),.d(in444),.sel(cs[1:0]),.out(muxpo12));
mux42 mux42p13(.a(in13),.b(in157),.c(in301),.d(in445),.sel(cs[1:0]),.out(muxpo13));
mux42 mux42p14(.a(in14),.b(in158),.c(in302),.d(in446),.sel(cs[1:0]),.out(muxpo14));
mux42 mux42p15(.a(in15),.b(in159),.c(in303),.d(in447),.sel(cs[1:0]),.out(muxpo15));
mux42 mux42p16(.a(in16),.b(in160),.c(in304),.d(in448),.sel(cs[1:0]),.out(muxpo16));
mux42 mux42p17(.a(in17),.b(in161),.c(in305),.d(in449),.sel(cs[1:0]),.out(muxpo17));
mux42 mux42p18(.a(in18),.b(in162),.c(in306),.d(in450),.sel(cs[1:0]),.out(muxpo18));
mux42 mux42p19(.a(in19),.b(in163),.c(in307),.d(in451),.sel(cs[1:0]),.out(muxpo19));
mux42 mux42p20(.a(in20),.b(in164),.c(in308),.d(in452),.sel(cs[1:0]),.out(muxpo20));
mux42 mux42p21(.a(in21),.b(in165),.c(in309),.d(in453),.sel(cs[1:0]),.out(muxpo21));
mux42 mux42p22(.a(in22),.b(in166),.c(in310),.d(in454),.sel(cs[1:0]),.out(muxpo22));
mux42 mux42p23(.a(in23),.b(in167),.c(in311),.d(in455),.sel(cs[1:0]),.out(muxpo23));
mux42 mux42p24(.a(in24),.b(in168),.c(in312),.d(in456),.sel(cs[1:0]),.out(muxpo24));
mux42 mux42p25(.a(in25),.b(in169),.c(in313),.d(in457),.sel(cs[1:0]),.out(muxpo25));
mux42 mux42p26(.a(in26),.b(in170),.c(in314),.d(in458),.sel(cs[1:0]),.out(muxpo26));
mux42 mux42p27(.a(in27),.b(in171),.c(in315),.d(in459),.sel(cs[1:0]),.out(muxpo27));
mux42 mux42p28(.a(in28),.b(in172),.c(in316),.d(in460),.sel(cs[1:0]),.out(muxpo28));
mux42 mux42p29(.a(in29),.b(in173),.c(in317),.d(in461),.sel(cs[1:0]),.out(muxpo29));
mux42 mux42p30(.a(in30),.b(in174),.c(in318),.d(in462),.sel(cs[1:0]),.out(muxpo30));
mux42 mux42p31(.a(in31),.b(in175),.c(in319),.d(in463),.sel(cs[1:0]),.out(muxpo31));
mux42 mux42p32(.a(in32),.b(in176),.c(in320),.d(in464),.sel(cs[1:0]),.out(muxpo32));
mux42 mux42p33(.a(in33),.b(in177),.c(in321),.d(in465),.sel(cs[1:0]),.out(muxpo33));
mux42 mux42p34(.a(in34),.b(in178),.c(in322),.d(in466),.sel(cs[1:0]),.out(muxpo34));
mux42 mux42p35(.a(in35),.b(in179),.c(in323),.d(in467),.sel(cs[1:0]),.out(muxpo35));
mux42 mux42p36(.a(in36),.b(in180),.c(in324),.d(in468),.sel(cs[1:0]),.out(muxpo36));
mux42 mux42p37(.a(in37),.b(in181),.c(in325),.d(in469),.sel(cs[1:0]),.out(muxpo37));
mux42 mux42p38(.a(in38),.b(in182),.c(in326),.d(in470),.sel(cs[1:0]),.out(muxpo38));
mux42 mux42p39(.a(in39),.b(in183),.c(in327),.d(in471),.sel(cs[1:0]),.out(muxpo39));
mux42 mux42p40(.a(in40),.b(in184),.c(in328),.d(in472),.sel(cs[1:0]),.out(muxpo40));
mux42 mux42p41(.a(in41),.b(in185),.c(in329),.d(in473),.sel(cs[1:0]),.out(muxpo41));
mux42 mux42p42(.a(in42),.b(in186),.c(in330),.d(in474),.sel(cs[1:0]),.out(muxpo42));
mux42 mux42p43(.a(in43),.b(in187),.c(in331),.d(in475),.sel(cs[1:0]),.out(muxpo43));
mux42 mux42p44(.a(in44),.b(in188),.c(in332),.d(in476),.sel(cs[1:0]),.out(muxpo44));
mux42 mux42p45(.a(in45),.b(in189),.c(in333),.d(in477),.sel(cs[1:0]),.out(muxpo45));
mux42 mux42p46(.a(in46),.b(in190),.c(in334),.d(in478),.sel(cs[1:0]),.out(muxpo46));
mux42 mux42p47(.a(in47),.b(in191),.c(in335),.d(in479),.sel(cs[1:0]),.out(muxpo47));
mux42 mux42p48(.a(in48),.b(in192),.c(in336),.d(in480),.sel(cs[1:0]),.out(muxpo48));
mux42 mux42p49(.a(in49),.b(in193),.c(in337),.d(in481),.sel(cs[1:0]),.out(muxpo49));
mux42 mux42p50(.a(in50),.b(in194),.c(in338),.d(in482),.sel(cs[1:0]),.out(muxpo50));
mux42 mux42p51(.a(in51),.b(in195),.c(in339),.d(in483),.sel(cs[1:0]),.out(muxpo51));
mux42 mux42p52(.a(in52),.b(in196),.c(in340),.d(in484),.sel(cs[1:0]),.out(muxpo52));
mux42 mux42p53(.a(in53),.b(in197),.c(in341),.d(in485),.sel(cs[1:0]),.out(muxpo53));
mux42 mux42p54(.a(in54),.b(in198),.c(in342),.d(in486),.sel(cs[1:0]),.out(muxpo54));
mux42 mux42p55(.a(in55),.b(in199),.c(in343),.d(in487),.sel(cs[1:0]),.out(muxpo55));
mux42 mux42p56(.a(in56),.b(in200),.c(in344),.d(in488),.sel(cs[1:0]),.out(muxpo56));
mux42 mux42p57(.a(in57),.b(in201),.c(in345),.d(in489),.sel(cs[1:0]),.out(muxpo57));
mux42 mux42p58(.a(in58),.b(in202),.c(in346),.d(in490),.sel(cs[1:0]),.out(muxpo58));
mux42 mux42p59(.a(in59),.b(in203),.c(in347),.d(in491),.sel(cs[1:0]),.out(muxpo59));
mux42 mux42p60(.a(in60),.b(in204),.c(in348),.d(in492),.sel(cs[1:0]),.out(muxpo60));
mux42 mux42p61(.a(in61),.b(in205),.c(in349),.d(in493),.sel(cs[1:0]),.out(muxpo61));
mux42 mux42p62(.a(in62),.b(in206),.c(in350),.d(in494),.sel(cs[1:0]),.out(muxpo62));
mux42 mux42p63(.a(in63),.b(in207),.c(in351),.d(in495),.sel(cs[1:0]),.out(muxpo63));
mux42 mux42p64(.a(in64),.b(in208),.c(in352),.d(in496),.sel(cs[1:0]),.out(muxpo64));
mux42 mux42p65(.a(in65),.b(in209),.c(in353),.d(in497),.sel(cs[1:0]),.out(muxpo65));
mux42 mux42p66(.a(in66),.b(in210),.c(in354),.d(in498),.sel(cs[1:0]),.out(muxpo66));
mux42 mux42p67(.a(in67),.b(in211),.c(in355),.d(in499),.sel(cs[1:0]),.out(muxpo67));
mux42 mux42p68(.a(in68),.b(in212),.c(in356),.d(in500),.sel(cs[1:0]),.out(muxpo68));
mux42 mux42p69(.a(in69),.b(in213),.c(in357),.d(in501),.sel(cs[1:0]),.out(muxpo69));
mux42 mux42p70(.a(in70),.b(in214),.c(in358),.d(in502),.sel(cs[1:0]),.out(muxpo70));
mux42 mux42p71(.a(in71),.b(in215),.c(in359),.d(in503),.sel(cs[1:0]),.out(muxpo71));
mux42 mux42p72(.a(in72),.b(in216),.c(in360),.d(in504),.sel(cs[1:0]),.out(muxpo72));
mux42 mux42p73(.a(in73),.b(in217),.c(in361),.d(in505),.sel(cs[1:0]),.out(muxpo73));
mux42 mux42p74(.a(in74),.b(in218),.c(in362),.d(in506),.sel(cs[1:0]),.out(muxpo74));
mux42 mux42p75(.a(in75),.b(in219),.c(in363),.d(in507),.sel(cs[1:0]),.out(muxpo75));
mux42 mux42p76(.a(in76),.b(in220),.c(in364),.d(in508),.sel(cs[1:0]),.out(muxpo76));
mux42 mux42p77(.a(in77),.b(in221),.c(in365),.d(in509),.sel(cs[1:0]),.out(muxpo77));
mux42 mux42p78(.a(in78),.b(in222),.c(in366),.d(in510),.sel(cs[1:0]),.out(muxpo78));
mux42 mux42p79(.a(in79),.b(in223),.c(in367),.d(in511),.sel(cs[1:0]),.out(muxpo79));
mux42 mux42p80(.a(in80),.b(in224),.c(in368),.d(in512),.sel(cs[1:0]),.out(muxpo80));
mux42 mux42p81(.a(in81),.b(in225),.c(in369),.d(in513),.sel(cs[1:0]),.out(muxpo81));
mux42 mux42p82(.a(in82),.b(in226),.c(in370),.d(in514),.sel(cs[1:0]),.out(muxpo82));
mux42 mux42p83(.a(in83),.b(in227),.c(in371),.d(in515),.sel(cs[1:0]),.out(muxpo83));
mux42 mux42p84(.a(in84),.b(in228),.c(in372),.d(in516),.sel(cs[1:0]),.out(muxpo84));
mux42 mux42p85(.a(in85),.b(in229),.c(in373),.d(in517),.sel(cs[1:0]),.out(muxpo85));
mux42 mux42p86(.a(in86),.b(in230),.c(in374),.d(in518),.sel(cs[1:0]),.out(muxpo86));
mux42 mux42p87(.a(in87),.b(in231),.c(in375),.d(in519),.sel(cs[1:0]),.out(muxpo87));
mux42 mux42p88(.a(in88),.b(in232),.c(in376),.d(in520),.sel(cs[1:0]),.out(muxpo88));
mux42 mux42p89(.a(in89),.b(in233),.c(in377),.d(in521),.sel(cs[1:0]),.out(muxpo89));
mux42 mux42p90(.a(in90),.b(in234),.c(in378),.d(in522),.sel(cs[1:0]),.out(muxpo90));
mux42 mux42p91(.a(in91),.b(in235),.c(in379),.d(in523),.sel(cs[1:0]),.out(muxpo91));
mux42 mux42p92(.a(in92),.b(in236),.c(in380),.d(in524),.sel(cs[1:0]),.out(muxpo92));
mux42 mux42p93(.a(in93),.b(in237),.c(in381),.d(in525),.sel(cs[1:0]),.out(muxpo93));
mux42 mux42p94(.a(in94),.b(in238),.c(in382),.d(in526),.sel(cs[1:0]),.out(muxpo94));
mux42 mux42p95(.a(in95),.b(in239),.c(in383),.d(in527),.sel(cs[1:0]),.out(muxpo95));
mux42 mux42p96(.a(in96),.b(in240),.c(in384),.d(in528),.sel(cs[1:0]),.out(muxpo96));
mux42 mux42p97(.a(in97),.b(in241),.c(in385),.d(in529),.sel(cs[1:0]),.out(muxpo97));
mux42 mux42p98(.a(in98),.b(in242),.c(in386),.d(in530),.sel(cs[1:0]),.out(muxpo98));
mux42 mux42p99(.a(in99),.b(in243),.c(in387),.d(in531),.sel(cs[1:0]),.out(muxpo99));
mux42 mux42p100(.a(in100),.b(in244),.c(in388),.d(in532),.sel(cs[1:0]),.out(muxpo100));
mux42 mux42p101(.a(in101),.b(in245),.c(in389),.d(in533),.sel(cs[1:0]),.out(muxpo101));
mux42 mux42p102(.a(in102),.b(in246),.c(in390),.d(in534),.sel(cs[1:0]),.out(muxpo102));
mux42 mux42p103(.a(in103),.b(in247),.c(in391),.d(in535),.sel(cs[1:0]),.out(muxpo103));
mux42 mux42p104(.a(in104),.b(in248),.c(in392),.d(in536),.sel(cs[1:0]),.out(muxpo104));
mux42 mux42p105(.a(in105),.b(in249),.c(in393),.d(in537),.sel(cs[1:0]),.out(muxpo105));
mux42 mux42p106(.a(in106),.b(in250),.c(in394),.d(in538),.sel(cs[1:0]),.out(muxpo106));
mux42 mux42p107(.a(in107),.b(in251),.c(in395),.d(in539),.sel(cs[1:0]),.out(muxpo107));
mux42 mux42p108(.a(in108),.b(in252),.c(in396),.d(in540),.sel(cs[1:0]),.out(muxpo108));
mux42 mux42p109(.a(in109),.b(in253),.c(in397),.d(in541),.sel(cs[1:0]),.out(muxpo109));
mux42 mux42p110(.a(in110),.b(in254),.c(in398),.d(in542),.sel(cs[1:0]),.out(muxpo110));
mux42 mux42p111(.a(in111),.b(in255),.c(in399),.d(in543),.sel(cs[1:0]),.out(muxpo111));
mux42 mux42p112(.a(in112),.b(in256),.c(in400),.d(in544),.sel(cs[1:0]),.out(muxpo112));
mux42 mux42p113(.a(in113),.b(in257),.c(in401),.d(in545),.sel(cs[1:0]),.out(muxpo113));
mux42 mux42p114(.a(in114),.b(in258),.c(in402),.d(in546),.sel(cs[1:0]),.out(muxpo114));
mux42 mux42p115(.a(in115),.b(in259),.c(in403),.d(in547),.sel(cs[1:0]),.out(muxpo115));
mux42 mux42p116(.a(in116),.b(in260),.c(in404),.d(in548),.sel(cs[1:0]),.out(muxpo116));
mux42 mux42p117(.a(in117),.b(in261),.c(in405),.d(in549),.sel(cs[1:0]),.out(muxpo117));
mux42 mux42p118(.a(in118),.b(in262),.c(in406),.d(in550),.sel(cs[1:0]),.out(muxpo118));
mux42 mux42p119(.a(in119),.b(in263),.c(in407),.d(in551),.sel(cs[1:0]),.out(muxpo119));
mux42 mux42p120(.a(in120),.b(in264),.c(in408),.d(in552),.sel(cs[1:0]),.out(muxpo120));
mux42 mux42p121(.a(in121),.b(in265),.c(in409),.d(in553),.sel(cs[1:0]),.out(muxpo121));
mux42 mux42p122(.a(in122),.b(in266),.c(in410),.d(in554),.sel(cs[1:0]),.out(muxpo122));
mux42 mux42p123(.a(in123),.b(in267),.c(in411),.d(in555),.sel(cs[1:0]),.out(muxpo123));
mux42 mux42p124(.a(in124),.b(in268),.c(in412),.d(in556),.sel(cs[1:0]),.out(muxpo124));
mux42 mux42p125(.a(in125),.b(in269),.c(in413),.d(in557),.sel(cs[1:0]),.out(muxpo125));
mux42 mux42p126(.a(in126),.b(in270),.c(in414),.d(in558),.sel(cs[1:0]),.out(muxpo126));
mux42 mux42p127(.a(in127),.b(in271),.c(in415),.d(in559),.sel(cs[1:0]),.out(muxpo127));
mux42 mux42p128(.a(in128),.b(in272),.c(in416),.d(in560),.sel(cs[1:0]),.out(muxpo128));
mux42 mux42p129(.a(in129),.b(in273),.c(in417),.d(in561),.sel(cs[1:0]),.out(muxpo129));
mux42 mux42p130(.a(in130),.b(in274),.c(in418),.d(in562),.sel(cs[1:0]),.out(muxpo130));
mux42 mux42p131(.a(in131),.b(in275),.c(in419),.d(in563),.sel(cs[1:0]),.out(muxpo131));
mux42 mux42p132(.a(in132),.b(in276),.c(in420),.d(in564),.sel(cs[1:0]),.out(muxpo132));
mux42 mux42p133(.a(in133),.b(in277),.c(in421),.d(in565),.sel(cs[1:0]),.out(muxpo133));
mux42 mux42p134(.a(in134),.b(in278),.c(in422),.d(in566),.sel(cs[1:0]),.out(muxpo134));
mux42 mux42p135(.a(in135),.b(in279),.c(in423),.d(in567),.sel(cs[1:0]),.out(muxpo135));
mux42 mux42p136(.a(in136),.b(in280),.c(in424),.d(in568),.sel(cs[1:0]),.out(muxpo136));
mux42 mux42p137(.a(in137),.b(in281),.c(in425),.d(in569),.sel(cs[1:0]),.out(muxpo137));
mux42 mux42p138(.a(in138),.b(in282),.c(in426),.d(in570),.sel(cs[1:0]),.out(muxpo138));
mux42 mux42p139(.a(in139),.b(in283),.c(in427),.d(in571),.sel(cs[1:0]),.out(muxpo139));
mux42 mux42p140(.a(in140),.b(in284),.c(in428),.d(in572),.sel(cs[1:0]),.out(muxpo140));
mux42 mux42p141(.a(in141),.b(in285),.c(in429),.d(in573),.sel(cs[1:0]),.out(muxpo141));
mux42 mux42p142(.a(in142),.b(in286),.c(in430),.d(in574),.sel(cs[1:0]),.out(muxpo142));
mux42 mux42p143(.a(in143),.b(in287),.c(in431),.d(in575),.sel(cs[1:0]),.out(muxpo143));



poolingfilter poolinfilter0(.in1(muxpo0),.in2(muxpo1),.in3(muxpo12),.in4(muxpo13),.out(muxpi0));
poolingfilter poolinfilter1(.in1(muxpo2),.in2(muxpo3),.in3(muxpo14),.in4(muxpo15),.out(muxpi1));
poolingfilter poolinfilter2(.in1(muxpo4),.in2(muxpo5),.in3(muxpo16),.in4(muxpo17),.out(muxpi2));
poolingfilter poolinfilter3(.in1(muxpo6),.in2(muxpo7),.in3(muxpo18),.in4(muxpo19),.out(muxpi3));
poolingfilter poolinfilter4(.in1(muxpo8),.in2(muxpo9),.in3(muxpo20),.in4(muxpo21),.out(muxpi4));
poolingfilter poolinfilter5(.in1(muxpo10),.in2(muxpo11),.in3(muxpo22),.in4(muxpo23),.out(muxpi5));
poolingfilter poolinfilter6(.in1(muxpo24),.in2(muxpo25),.in3(muxpo36),.in4(muxpo37),.out(muxpi6));
poolingfilter poolinfilter7(.in1(muxpo26),.in2(muxpo27),.in3(muxpo38),.in4(muxpo39),.out(muxpi7));
poolingfilter poolinfilter8(.in1(muxpo28),.in2(muxpo29),.in3(muxpo40),.in4(muxpo41),.out(muxpi8));
poolingfilter poolinfilter9(.in1(muxpo30),.in2(muxpo31),.in3(muxpo42),.in4(muxpo43),.out(muxpi9));
poolingfilter poolinfilter10(.in1(muxpo32),.in2(muxpo33),.in3(muxpo44),.in4(muxpo45),.out(muxpi10));
poolingfilter poolinfilter11(.in1(muxpo34),.in2(muxpo35),.in3(muxpo46),.in4(muxpo47),.out(muxpi11));
poolingfilter poolinfilter12(.in1(muxpo48),.in2(muxpo49),.in3(muxpo60),.in4(muxpo61),.out(muxpi12));
poolingfilter poolinfilter13(.in1(muxpo50),.in2(muxpo51),.in3(muxpo62),.in4(muxpo63),.out(muxpi13));
poolingfilter poolinfilter14(.in1(muxpo52),.in2(muxpo53),.in3(muxpo64),.in4(muxpo65),.out(muxpi14));
poolingfilter poolinfilter15(.in1(muxpo54),.in2(muxpo55),.in3(muxpo66),.in4(muxpo67),.out(muxpi15));
poolingfilter poolinfilter16(.in1(muxpo56),.in2(muxpo57),.in3(muxpo68),.in4(muxpo69),.out(muxpi16));
poolingfilter poolinfilter17(.in1(muxpo58),.in2(muxpo59),.in3(muxpo70),.in4(muxpo71),.out(muxpi17));
poolingfilter poolinfilter18(.in1(muxpo72),.in2(muxpo73),.in3(muxpo84),.in4(muxpo85),.out(muxpi18));
poolingfilter poolinfilter19(.in1(muxpo74),.in2(muxpo75),.in3(muxpo86),.in4(muxpo87),.out(muxpi19));
poolingfilter poolinfilter20(.in1(muxpo76),.in2(muxpo77),.in3(muxpo88),.in4(muxpo89),.out(muxpi20));
poolingfilter poolinfilter21(.in1(muxpo78),.in2(muxpo79),.in3(muxpo90),.in4(muxpo91),.out(muxpi21));
poolingfilter poolinfilter22(.in1(muxpo80),.in2(muxpo81),.in3(muxpo92),.in4(muxpo93),.out(muxpi22));
poolingfilter poolinfilter23(.in1(muxpo82),.in2(muxpo83),.in3(muxpo94),.in4(muxpo95),.out(muxpi23));
poolingfilter poolinfilter24(.in1(muxpo96),.in2(muxpo97),.in3(muxpo108),.in4(muxpo109),.out(muxpi24));
poolingfilter poolinfilter25(.in1(muxpo98),.in2(muxpo99),.in3(muxpo110),.in4(muxpo111),.out(muxpi25));
poolingfilter poolinfilter26(.in1(muxpo100),.in2(muxpo101),.in3(muxpo112),.in4(muxpo113),.out(muxpi26));
poolingfilter poolinfilter27(.in1(muxpo102),.in2(muxpo103),.in3(muxpo114),.in4(muxpo115),.out(muxpi27));
poolingfilter poolinfilter28(.in1(muxpo104),.in2(muxpo105),.in3(muxpo116),.in4(muxpo117),.out(muxpi28));
poolingfilter poolinfilter29(.in1(muxpo106),.in2(muxpo107),.in3(muxpo118),.in4(muxpo119),.out(muxpi29));
poolingfilter poolinfilter30(.in1(muxpo120),.in2(muxpo121),.in3(muxpo132),.in4(muxpo133),.out(muxpi30));
poolingfilter poolinfilter31(.in1(muxpo122),.in2(muxpo123),.in3(muxpo134),.in4(muxpo135),.out(muxpi31));
poolingfilter poolinfilter32(.in1(muxpo124),.in2(muxpo125),.in3(muxpo136),.in4(muxpo137),.out(muxpi32));
poolingfilter poolinfilter33(.in1(muxpo126),.in2(muxpo127),.in3(muxpo138),.in4(muxpo139),.out(muxpi33));
poolingfilter poolinfilter34(.in1(muxpo128),.in2(muxpo129),.in3(muxpo140),.in4(muxpo141),.out(muxpi34));
poolingfilter poolinfilter35(.in1(muxpo130),.in2(muxpo131),.in3(muxpo142),.in4(muxpo143),.out(muxpi35));


/*
demux42 demuxp0(.a(out0),.b(out36),.c(out72),.d(out108),.sel(cs[1:0]),.out(muxpi0));
demux42 demuxp1(.a(out1),.b(out37),.c(out73),.d(out109),.sel(cs[1:0]),.out(muxpi1));
demux42 demuxp2(.a(out2),.b(out38),.c(out74),.d(out110),.sel(cs[1:0]),.out(muxpi2));
demux42 demuxp3(.a(out3),.b(out39),.c(out75),.d(out111),.sel(cs[1:0]),.out(muxpi3));
demux42 demuxp4(.a(out4),.b(out40),.c(out76),.d(out112),.sel(cs[1:0]),.out(muxpi4));
demux42 demuxp5(.a(out5),.b(out41),.c(out77),.d(out113),.sel(cs[1:0]),.out(muxpi5));
demux42 demuxp6(.a(out6),.b(out42),.c(out78),.d(out114),.sel(cs[1:0]),.out(muxpi6));
demux42 demuxp7(.a(out7),.b(out43),.c(out79),.d(out115),.sel(cs[1:0]),.out(muxpi7));
demux42 demuxp8(.a(out8),.b(out44),.c(out80),.d(out116),.sel(cs[1:0]),.out(muxpi8));
demux42 demuxp9(.a(out9),.b(out45),.c(out81),.d(out117),.sel(cs[1:0]),.out(muxpi9));
demux42 demuxp10(.a(out10),.b(out46),.c(out82),.d(out118),.sel(cs[1:0]),.out(muxpi10));
demux42 demuxp11(.a(out11),.b(out47),.c(out83),.d(out119),.sel(cs[1:0]),.out(muxpi11));
demux42 demuxp12(.a(out12),.b(out48),.c(out84),.d(out120),.sel(cs[1:0]),.out(muxpi12));
demux42 demuxp13(.a(out13),.b(out49),.c(out85),.d(out121),.sel(cs[1:0]),.out(muxpi13));
demux42 demuxp14(.a(out14),.b(out50),.c(out86),.d(out122),.sel(cs[1:0]),.out(muxpi14));
demux42 demuxp15(.a(out15),.b(out51),.c(out87),.d(out123),.sel(cs[1:0]),.out(muxpi15));
demux42 demuxp16(.a(out16),.b(out52),.c(out88),.d(out124),.sel(cs[1:0]),.out(muxpi16));
demux42 demuxp17(.a(out17),.b(out53),.c(out89),.d(out125),.sel(cs[1:0]),.out(muxpi17));
demux42 demuxp18(.a(out18),.b(out54),.c(out90),.d(out126),.sel(cs[1:0]),.out(muxpi18));
demux42 demuxp19(.a(out19),.b(out55),.c(out91),.d(out127),.sel(cs[1:0]),.out(muxpi19));
demux42 demuxp20(.a(out20),.b(out56),.c(out92),.d(out128),.sel(cs[1:0]),.out(muxpi20));
demux42 demuxp21(.a(out21),.b(out57),.c(out93),.d(out129),.sel(cs[1:0]),.out(muxpi21));
demux42 demuxp22(.a(out22),.b(out58),.c(out94),.d(out130),.sel(cs[1:0]),.out(muxpi22));
demux42 demuxp23(.a(out23),.b(out59),.c(out95),.d(out131),.sel(cs[1:0]),.out(muxpi23));
demux42 demuxp24(.a(out24),.b(out60),.c(out96),.d(out132),.sel(cs[1:0]),.out(muxpi24));
demux42 demuxp25(.a(out25),.b(out61),.c(out97),.d(out133),.sel(cs[1:0]),.out(muxpi25));
demux42 demuxp26(.a(out26),.b(out62),.c(out98),.d(out134),.sel(cs[1:0]),.out(muxpi26));
demux42 demuxp27(.a(out27),.b(out63),.c(out99),.d(out135),.sel(cs[1:0]),.out(muxpi27));
demux42 demuxp28(.a(out28),.b(out64),.c(out100),.d(out136),.sel(cs[1:0]),.out(muxpi28));
demux42 demuxp29(.a(out29),.b(out65),.c(out101),.d(out137),.sel(cs[1:0]),.out(muxpi29));
demux42 demuxp30(.a(out30),.b(out66),.c(out102),.d(out138),.sel(cs[1:0]),.out(muxpi30));
demux42 demuxp31(.a(out31),.b(out67),.c(out103),.d(out139),.sel(cs[1:0]),.out(muxpi31));
demux42 demuxp32(.a(out32),.b(out68),.c(out104),.d(out140),.sel(cs[1:0]),.out(muxpi32));
demux42 demuxp33(.a(out33),.b(out69),.c(out105),.d(out141),.sel(cs[1:0]),.out(muxpi33));
demux42 demuxp34(.a(out34),.b(out70),.c(out106),.d(out142),.sel(cs[1:0]),.out(muxpi34));
demux42 demuxp35(.a(out35),.b(out71),.c(out107),.d(out143),.sel(cs[1:0]),.out(muxpi35));
*/

localparam WAIT = 3'b000;
localparam CALC1 = 3'b001;
localparam CALC2 = 3'b010;
localparam CALC3 = 3'b011;
localparam CALC4 = 3'b100;
localparam READY = 3'b101;
localparam START = 3'b111;

reg ready;
reg [2:0] state;
reg [2:0] next_state;
reg [2:0] cs;



always @(posedge clk or posedge start)
	begin
	if (start)begin
	next_state <= START;
	ready <= 0;
	end
	else
	begin
	state <= next_state;
	end
	case(state)
		START:
		begin
			next_state <= CALC1;
			cs <= 3'b000;
		end
		CALC1:
		begin
			muxreg0<=muxpi0;muxreg1<=muxpi1;muxreg2<=muxpi2;muxreg3<=muxpi3;muxreg4<=muxpi4;muxreg5<=muxpi5;muxreg6<=muxpi6;muxreg7<=muxpi7;muxreg8<=muxpi8;muxreg9<=muxpi9;muxreg10<=muxpi10;muxreg11<=muxpi11;muxreg12<=muxpi12;muxreg13<=muxpi13;muxreg14<=muxpi14;muxreg15<=muxpi15;muxreg16<=muxpi16;muxreg17<=muxpi17;muxreg18<=muxpi18;muxreg19<=muxpi19;muxreg20<=muxpi20;muxreg21<=muxpi21;muxreg22<=muxpi22;muxreg23<=muxpi23;muxreg24<=muxpi24;muxreg25<=muxpi25;muxreg26<=muxpi26;muxreg27<=muxpi27;muxreg28<=muxpi28;muxreg29<=muxpi29;muxreg30<=muxpi30;muxreg31<=muxpi31;muxreg32<=muxpi32;muxreg33<=muxpi33;muxreg34<=muxpi34;muxreg35<=muxpi35;
			next_state <= CALC2;
			cs <= 3'b000;
		end
		CALC2:
		begin
			muxreg36<=muxpi0;muxreg37<=muxpi1;muxreg38<=muxpi2;muxreg39<=muxpi3;muxreg40<=muxpi4;muxreg41<=muxpi5;muxreg42<=muxpi6;muxreg43<=muxpi7;muxreg44<=muxpi8;muxreg45<=muxpi9;muxreg46<=muxpi10;muxreg47<=muxpi11;muxreg48<=muxpi12;muxreg49<=muxpi13;muxreg50<=muxpi14;muxreg51<=muxpi15;muxreg52<=muxpi16;muxreg53<=muxpi17;muxreg54<=muxpi18;muxreg55<=muxpi19;muxreg56<=muxpi20;muxreg57<=muxpi21;muxreg58<=muxpi22;muxreg59<=muxpi23;muxreg60<=muxpi24;muxreg61<=muxpi25;muxreg62<=muxpi26;muxreg63<=muxpi27;muxreg64<=muxpi28;muxreg65<=muxpi29;muxreg66<=muxpi30;muxreg67<=muxpi31;muxreg68<=muxpi32;muxreg69<=muxpi33;muxreg70<=muxpi34;muxreg71<=muxpi35;
			next_state <= CALC3;
			cs <= 3'b001;
		end
		CALC3:
		begin
			muxreg72<=muxpi0;muxreg73<=muxpi1;muxreg74<=muxpi2;muxreg75<=muxpi3;muxreg76<=muxpi4;muxreg77<=muxpi5;muxreg78<=muxpi6;muxreg79<=muxpi7;muxreg80<=muxpi8;muxreg81<=muxpi9;muxreg82<=muxpi10;muxreg83<=muxpi11;muxreg84<=muxpi12;muxreg85<=muxpi13;muxreg86<=muxpi14;muxreg87<=muxpi15;muxreg88<=muxpi16;muxreg89<=muxpi17;muxreg90<=muxpi18;muxreg91<=muxpi19;muxreg92<=muxpi20;muxreg93<=muxpi21;muxreg94<=muxpi22;muxreg95<=muxpi23;muxreg96<=muxpi24;muxreg97<=muxpi25;muxreg98<=muxpi26;muxreg99<=muxpi27;muxreg100<=muxpi28;muxreg101<=muxpi29;muxreg102<=muxpi30;muxreg103<=muxpi31;muxreg104<=muxpi32;muxreg105<=muxpi33;muxreg106<=muxpi34;muxreg107<=muxpi35;
			next_state <= CALC4;
			cs <= 3'b010;
		end
		CALC4:
		begin
			 muxreg108<=muxpi0;muxreg109<=muxpi1;muxreg110<=muxpi2;muxreg111<=muxpi3;muxreg112<=muxpi4;muxreg113<=muxpi5;muxreg114<=muxpi6;muxreg115<=muxpi7;muxreg116<=muxpi8;muxreg117<=muxpi9;muxreg118<=muxpi10;muxreg119<=muxpi11;muxreg120<=muxpi12;muxreg121<=muxpi13;muxreg122<=muxpi14;muxreg123<=muxpi15;muxreg124<=muxpi16;muxreg125<=muxpi17;muxreg126<=muxpi18;muxreg127<=muxpi19;muxreg128<=muxpi20;muxreg129<=muxpi21;muxreg130<=muxpi22;muxreg131<=muxpi23;muxreg132<=muxpi24;muxreg133<=muxpi25;muxreg134<=muxpi26;muxreg135<=muxpi27;muxreg136<=muxpi28;muxreg137<=muxpi29;muxreg138<=muxpi30;muxreg139<=muxpi31;muxreg140<=muxpi32;muxreg141<=muxpi33;muxreg142<=muxpi34;muxreg143<=muxpi35;
			next_state <= READY;
			cs <= 3'b011;
			ready <= 1;
		end
		READY:
		begin
			next_state <= WAIT;
			cs <= 3'b100;
			ready <= 0;
		end
		/*default:
		begin
			state <= WAIT;
			cs <= 3'b000;
		end*/
		endcase
	end
	
	 assign out0=muxreg0;assign out1=muxreg1;assign out2=muxreg2;assign out3=muxreg3;assign out4=muxreg4;assign out5=muxreg5;assign out6=muxreg6;assign out7=muxreg7;assign out8=muxreg8;assign out9=muxreg9;assign out10=muxreg10;assign out11=muxreg11;assign out12=muxreg12;assign out13=muxreg13;assign out14=muxreg14;assign out15=muxreg15;assign out16=muxreg16;assign out17=muxreg17;assign out18=muxreg18;assign out19=muxreg19;assign out20=muxreg20;assign out21=muxreg21;assign out22=muxreg22;assign out23=muxreg23;assign out24=muxreg24;assign out25=muxreg25;assign out26=muxreg26;assign out27=muxreg27;assign out28=muxreg28;assign out29=muxreg29;assign out30=muxreg30;assign out31=muxreg31;assign out32=muxreg32;assign out33=muxreg33;assign out34=muxreg34;assign out35=muxreg35;assign out36=muxreg36;assign out37=muxreg37;assign out38=muxreg38;assign out39=muxreg39;assign out40=muxreg40;assign out41=muxreg41;assign out42=muxreg42;assign out43=muxreg43;assign out44=muxreg44;assign out45=muxreg45;assign out46=muxreg46;assign out47=muxreg47;assign out48=muxreg48;assign out49=muxreg49;assign out50=muxreg50;assign out51=muxreg51;assign out52=muxreg52;assign out53=muxreg53;assign out54=muxreg54;assign out55=muxreg55;assign out56=muxreg56;assign out57=muxreg57;assign out58=muxreg58;assign out59=muxreg59;assign out60=muxreg60;assign out61=muxreg61;assign out62=muxreg62;assign out63=muxreg63;assign out64=muxreg64;assign out65=muxreg65;assign out66=muxreg66;assign out67=muxreg67;assign out68=muxreg68;assign out69=muxreg69;assign out70=muxreg70;assign out71=muxreg71;assign out72=muxreg72;assign out73=muxreg73;assign out74=muxreg74;assign out75=muxreg75;assign out76=muxreg76;assign out77=muxreg77;assign out78=muxreg78;assign out79=muxreg79;assign out80=muxreg80;assign out81=muxreg81;assign out82=muxreg82;assign out83=muxreg83;assign out84=muxreg84;assign out85=muxreg85;assign out86=muxreg86;assign out87=muxreg87;assign out88=muxreg88;assign out89=muxreg89;assign out90=muxreg90;assign out91=muxreg91;assign out92=muxreg92;assign out93=muxreg93;assign out94=muxreg94;assign out95=muxreg95;assign out96=muxreg96;assign out97=muxreg97;assign out98=muxreg98;assign out99=muxreg99;assign out100=muxreg100;assign out101=muxreg101;assign out102=muxreg102;assign out103=muxreg103;assign out104=muxreg104;assign out105=muxreg105;assign out106=muxreg106;assign out107=muxreg107;assign out108=muxreg108;assign out109=muxreg109;assign out110=muxreg110;assign out111=muxreg111;assign out112=muxreg112;assign out113=muxreg113;assign out114=muxreg114;assign out115=muxreg115;assign out116=muxreg116;assign out117=muxreg117;assign out118=muxreg118;assign out119=muxreg119;assign out120=muxreg120;assign out121=muxreg121;assign out122=muxreg122;assign out123=muxreg123;assign out124=muxreg124;assign out125=muxreg125;assign out126=muxreg126;assign out127=muxreg127;assign out128=muxreg128;assign out129=muxreg129;assign out130=muxreg130;assign out131=muxreg131;assign out132=muxreg132;assign out133=muxreg133;assign out134=muxreg134;assign out135=muxreg135;assign out136=muxreg136;assign out137=muxreg137;assign out138=muxreg138;assign out139=muxreg139;assign out140=muxreg140;assign out141=muxreg141;assign out142=muxreg142;assign out143=muxreg143;

endmodule


