`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    00:44:38 11/03/2017 
// Design Name: 
// Module Name:    ConvLayer 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ConvLayer(weight0, weight1, weight2, weight3, weight4, weight5, weight6, weight7, 
weight8, weight9, weight10, weight11, weight12, weight13, weight14, weight15, weight16, 
weight17, weight18, weight19, weight20, weight21, weight22, weight23, weight24,in0,in1,in2,in3,in4,in5,in6,in7,in8,in9,in10,in11,in12,in13,in14,in15,in16,in17,in18,in19,in20,in21,in22,in23,in24,in25,in26,in27,in28,in29,in30,in31,in32,in33,in34,in35,in36,in37,in38,in39,in40,in41,in42,in43,in44,in45,in46,in47,in48,in49,in50,in51,in52,in53,in54,in55,in56,in57,in58,in59,in60,in61,in62,in63,in64,in65,in66,in67,in68,in69,in70,in71,in72,in73,in74,in75,in76,in77,in78,in79,in80,in81,in82,in83,in84,in85,in86,in87,in88,in89,in90,in91,in92,in93,in94,in95,in96,in97,in98,in99,in100,in101,in102,in103,in104,in105,in106,in107,in108,in109,in110,in111,in112,in113,in114,in115,in116,in117,in118,in119,in120,in121,in122,in123,in124,in125,in126,in127,in128,in129,in130,in131,in132,in133,in134,in135,in136,in137,in138,in139,in140,in141,in142,in143,in144,in145,in146,in147,in148,in149,in150,in151,in152,in153,in154,in155,in156,in157,in158,in159,in160,in161,in162,in163,in164,in165,in166,in167,in168,in169,in170,in171,in172,in173,in174,in175,in176,in177,in178,in179,in180,in181,in182,in183,in184,in185,in186,in187,in188,in189,in190,in191,in192,in193,in194,in195,in196,in197,in198,in199,in200,in201,in202,in203,in204,in205,in206,in207,in208,in209,in210,in211,in212,in213,in214,in215,in216,in217,in218,in219,in220,in221,in222,in223,in224,in225,in226,in227,in228,in229,in230,in231,in232,in233,in234,in235,in236,in237,in238,in239,in240,in241,in242,in243,in244,in245,in246,in247,in248,in249,in250,in251,in252,in253,in254,in255,in256,in257,in258,in259,in260,in261,in262,in263,in264,in265,in266,in267,in268,in269,in270,in271,in272,in273,in274,in275,in276,in277,in278,in279,in280,in281,in282,in283,in284,in285,in286,in287,in288,in289,in290,in291,in292,in293,in294,in295,in296,in297,in298,in299,in300,in301,in302,in303,in304,in305,in306,in307,in308,in309,in310,in311,in312,in313,in314,in315,in316,in317,in318,in319,in320,in321,in322,in323,in324,in325,in326,in327,in328,in329,in330,in331,in332,in333,in334,in335,in336,in337,in338,in339,in340,in341,in342,in343,in344,in345,in346,in347,in348,in349,in350,in351,in352,in353,in354,in355,in356,in357,in358,in359,in360,in361,in362,in363,in364,in365,in366,in367,in368,in369,in370,in371,in372,in373,in374,in375,in376,in377,in378,in379,in380,in381,in382,in383,in384,in385,in386,in387,in388,in389,in390,in391,in392,in393,in394,in395,in396,in397,in398,in399,in400,in401,in402,in403,in404,in405,in406,in407,in408,in409,in410,in411,in412,in413,in414,in415,in416,in417,in418,in419,in420,in421,in422,in423,in424,in425,in426,in427,in428,in429,in430,in431,in432,in433,in434,in435,in436,in437,in438,in439,in440,in441,in442,in443,in444,in445,in446,in447,in448,in449,in450,in451,in452,in453,in454,in455,in456,in457,in458,in459,in460,in461,in462,in463,in464,in465,in466,in467,in468,in469,in470,in471,in472,in473,in474,in475,in476,in477,in478,in479,in480,in481,in482,in483,in484,in485,in486,in487,in488,in489,in490,in491,in492,in493,in494,in495,in496,in497,in498,in499,in500,in501,in502,in503,in504,in505,in506,in507,in508,in509,in510,in511,in512,in513,in514,in515,in516,in517,in518,in519,in520,in521,in522,in523,in524,in525,in526,in527,in528,in529,in530,in531,in532,in533,in534,in535,in536,in537,in538,in539,in540,in541,in542,in543,in544,in545,in546,in547,in548,in549,in550,in551,in552,in553,in554,in555,in556,in557,in558,in559,in560,in561,in562,in563,in564,in565,in566,in567,in568,in569,in570,in571,in572,in573,in574,in575,in576,in577,in578,in579,in580,in581,in582,in583,in584,in585,in586,in587,in588,in589,in590,in591,in592,in593,in594,in595,in596,in597,in598,in599,in600,in601,in602,in603,in604,in605,in606,in607,in608,in609,in610,in611,in612,in613,in614,in615,in616,in617,in618,in619,in620,in621,in622,in623,in624,in625,in626,in627,in628,in629,in630,in631,in632,in633,in634,in635,in636,in637,in638,in639,in640,in641,in642,in643,in644,in645,in646,in647,in648,in649,in650,in651,in652,in653,in654,in655,in656,in657,in658,in659,in660,in661,in662,in663,in664,in665,in666,in667,in668,in669,in670,in671,in672,in673,in674,in675,in676,in677,in678,in679,in680,in681,in682,in683,in684,in685,in686,in687,in688,in689,in690,in691,in692,in693,in694,in695,in696,in697,in698,in699,in700,in701,in702,in703,in704,in705,in706,in707,in708,in709,in710,in711,in712,in713,in714,in715,in716,in717,in718,in719,in720,in721,in722,in723,in724,in725,in726,in727,in728,in729,in730,in731,in732,in733,in734,in735,in736,in737,in738,in739,in740,in741,in742,in743,in744,in745,in746,in747,in748,in749,in750,in751,in752,in753,in754,in755,in756,in757,in758,in759,in760,in761,in762,in763,in764,in765,in766,in767,in768,in769,in770,in771,in772,in773,in774,in775,in776,in777,in778,in779,in780,in781,in782,in783,
bias, clk,conv0,conv1,conv2,conv3,conv4,conv5,conv6,conv7,conv8,conv9,conv10,conv11,conv12,conv13,conv14,conv15,conv16,conv17,conv18,conv19,conv20,conv21,conv22,conv23,conv24,conv25,conv26,conv27,conv28,conv29,conv30,conv31,conv32,conv33,conv34,conv35,conv36,conv37,conv38,conv39,conv40,conv41,conv42,conv43,conv44,conv45,conv46,conv47,conv48,conv49,conv50,conv51,conv52,conv53,conv54,conv55,conv56,conv57,conv58,conv59,conv60,conv61,conv62,conv63,conv64,conv65,conv66,conv67,conv68,conv69,conv70,conv71,conv72,conv73,conv74,conv75,conv76,conv77,conv78,conv79,conv80,conv81,conv82,conv83,conv84,conv85,conv86,conv87,conv88,conv89,conv90,conv91,conv92,conv93,conv94,conv95,conv96,conv97,conv98,conv99,conv100,conv101,conv102,conv103,conv104,conv105,conv106,conv107,conv108,conv109,conv110,conv111,conv112,conv113,conv114,conv115,conv116,conv117,conv118,conv119,conv120,conv121,conv122,conv123,conv124,conv125,conv126,conv127,conv128,conv129,conv130,conv131,conv132,conv133,conv134,conv135,conv136,conv137,conv138,conv139,conv140,conv141,conv142,conv143,conv144,conv145,conv146,conv147,conv148,conv149,conv150,conv151,conv152,conv153,conv154,conv155,conv156,conv157,conv158,conv159,conv160,conv161,conv162,conv163,conv164,conv165,conv166,conv167,conv168,conv169,conv170,conv171,conv172,conv173,conv174,conv175,conv176,conv177,conv178,conv179,conv180,conv181,conv182,conv183,conv184,conv185,conv186,conv187,conv188,conv189,conv190,conv191,conv192,conv193,conv194,conv195,conv196,conv197,conv198,conv199,conv200,conv201,conv202,conv203,conv204,conv205,conv206,conv207,conv208,conv209,conv210,conv211,conv212,conv213,conv214,conv215,conv216,conv217,conv218,conv219,conv220,conv221,conv222,conv223,conv224,conv225,conv226,conv227,conv228,conv229,conv230,conv231,conv232,conv233,conv234,conv235,conv236,conv237,conv238,conv239,conv240,conv241,conv242,conv243,conv244,conv245,conv246,conv247,conv248,conv249,conv250,conv251,conv252,conv253,conv254,conv255,conv256,conv257,conv258,conv259,conv260,conv261,conv262,conv263,conv264,conv265,conv266,conv267,conv268,conv269,conv270,conv271,conv272,conv273,conv274,conv275,conv276,conv277,conv278,conv279,conv280,conv281,conv282,conv283,conv284,conv285,conv286,conv287,conv288,conv289,conv290,conv291,conv292,conv293,conv294,conv295,conv296,conv297,conv298,conv299,conv300,conv301,conv302,conv303,conv304,conv305,conv306,conv307,conv308,conv309,conv310,conv311,conv312,conv313,conv314,conv315,conv316,conv317,conv318,conv319,conv320,conv321,conv322,conv323,conv324,conv325,conv326,conv327,conv328,conv329,conv330,conv331,conv332,conv333,conv334,conv335,conv336,conv337,conv338,conv339,conv340,conv341,conv342,conv343,conv344,conv345,conv346,conv347,conv348,conv349,conv350,conv351,conv352,conv353,conv354,conv355,conv356,conv357,conv358,conv359,conv360,conv361,conv362,conv363,conv364,conv365,conv366,conv367,conv368,conv369,conv370,conv371,conv372,conv373,conv374,conv375,conv376,conv377,conv378,conv379,conv380,conv381,conv382,conv383,conv384,conv385,conv386,conv387,conv388,conv389,conv390,conv391,conv392,conv393,conv394,conv395,conv396,conv397,conv398,conv399,conv400,conv401,conv402,conv403,conv404,conv405,conv406,conv407,conv408,conv409,conv410,conv411,conv412,conv413,conv414,conv415,conv416,conv417,conv418,conv419,conv420,conv421,conv422,conv423,conv424,conv425,conv426,conv427,conv428,conv429,conv430,conv431,conv432,conv433,conv434,conv435,conv436,conv437,conv438,conv439,conv440,conv441,conv442,conv443,conv444,conv445,conv446,conv447,conv448,conv449,conv450,conv451,conv452,conv453,conv454,conv455,conv456,conv457,conv458,conv459,conv460,conv461,conv462,conv463,conv464,conv465,conv466,conv467,conv468,conv469,conv470,conv471,conv472,conv473,conv474,conv475,conv476,conv477,conv478,conv479,conv480,conv481,conv482,conv483,conv484,conv485,conv486,conv487,conv488,conv489,conv490,conv491,conv492,conv493,conv494,conv495,conv496,conv497,conv498,conv499,conv500,conv501,conv502,conv503,conv504,conv505,conv506,conv507,conv508,conv509,conv510,conv511,conv512,conv513,conv514,conv515,conv516,conv517,conv518,conv519,conv520,conv521,conv522,conv523,conv524,conv525,conv526,conv527,conv528,conv529,conv530,conv531,conv532,conv533,conv534,conv535,conv536,conv537,conv538,conv539,conv540,conv541,conv542,conv543,conv544,conv545,conv546,conv547,conv548,conv549,conv550,conv551,conv552,conv553,conv554,conv555,conv556,conv557,conv558,conv559,conv560,conv561,conv562,conv563,conv564,conv565,conv566,conv567,conv568,conv569,conv570,conv571,conv572,conv573,conv574,conv575,
ready,start);
	 
output ready;
reg ready;
input start;
input [7:0] in0;
input [7:0] in1;
input [7:0] in2;
input [7:0] in3;
input [7:0] in4;
input [7:0] in5;
input [7:0] in6;
input [7:0] in7;
input [7:0] in8;
input [7:0] in9;
input [7:0] in10;
input [7:0] in11;
input [7:0] in12;
input [7:0] in13;
input [7:0] in14;
input [7:0] in15;
input [7:0] in16;
input [7:0] in17;
input [7:0] in18;
input [7:0] in19;
input [7:0] in20;
input [7:0] in21;
input [7:0] in22;
input [7:0] in23;
input [7:0] in24;
input [7:0] in25;
input [7:0] in26;
input [7:0] in27;
input [7:0] in28;
input [7:0] in29;
input [7:0] in30;
input [7:0] in31;
input [7:0] in32;
input [7:0] in33;
input [7:0] in34;
input [7:0] in35;
input [7:0] in36;
input [7:0] in37;
input [7:0] in38;
input [7:0] in39;
input [7:0] in40;
input [7:0] in41;
input [7:0] in42;
input [7:0] in43;
input [7:0] in44;
input [7:0] in45;
input [7:0] in46;
input [7:0] in47;
input [7:0] in48;
input [7:0] in49;
input [7:0] in50;
input [7:0] in51;
input [7:0] in52;
input [7:0] in53;
input [7:0] in54;
input [7:0] in55;
input [7:0] in56;
input [7:0] in57;
input [7:0] in58;
input [7:0] in59;
input [7:0] in60;
input [7:0] in61;
input [7:0] in62;
input [7:0] in63;
input [7:0] in64;
input [7:0] in65;
input [7:0] in66;
input [7:0] in67;
input [7:0] in68;
input [7:0] in69;
input [7:0] in70;
input [7:0] in71;
input [7:0] in72;
input [7:0] in73;
input [7:0] in74;
input [7:0] in75;
input [7:0] in76;
input [7:0] in77;
input [7:0] in78;
input [7:0] in79;
input [7:0] in80;
input [7:0] in81;
input [7:0] in82;
input [7:0] in83;
input [7:0] in84;
input [7:0] in85;
input [7:0] in86;
input [7:0] in87;
input [7:0] in88;
input [7:0] in89;
input [7:0] in90;
input [7:0] in91;
input [7:0] in92;
input [7:0] in93;
input [7:0] in94;
input [7:0] in95;
input [7:0] in96;
input [7:0] in97;
input [7:0] in98;
input [7:0] in99;
input [7:0] in100;
input [7:0] in101;
input [7:0] in102;
input [7:0] in103;
input [7:0] in104;
input [7:0] in105;
input [7:0] in106;
input [7:0] in107;
input [7:0] in108;
input [7:0] in109;
input [7:0] in110;
input [7:0] in111;
input [7:0] in112;
input [7:0] in113;
input [7:0] in114;
input [7:0] in115;
input [7:0] in116;
input [7:0] in117;
input [7:0] in118;
input [7:0] in119;
input [7:0] in120;
input [7:0] in121;
input [7:0] in122;
input [7:0] in123;
input [7:0] in124;
input [7:0] in125;
input [7:0] in126;
input [7:0] in127;
input [7:0] in128;
input [7:0] in129;
input [7:0] in130;
input [7:0] in131;
input [7:0] in132;
input [7:0] in133;
input [7:0] in134;
input [7:0] in135;
input [7:0] in136;
input [7:0] in137;
input [7:0] in138;
input [7:0] in139;
input [7:0] in140;
input [7:0] in141;
input [7:0] in142;
input [7:0] in143;
input [7:0] in144;
input [7:0] in145;
input [7:0] in146;
input [7:0] in147;
input [7:0] in148;
input [7:0] in149;
input [7:0] in150;
input [7:0] in151;
input [7:0] in152;
input [7:0] in153;
input [7:0] in154;
input [7:0] in155;
input [7:0] in156;
input [7:0] in157;
input [7:0] in158;
input [7:0] in159;
input [7:0] in160;
input [7:0] in161;
input [7:0] in162;
input [7:0] in163;
input [7:0] in164;
input [7:0] in165;
input [7:0] in166;
input [7:0] in167;
input [7:0] in168;
input [7:0] in169;
input [7:0] in170;
input [7:0] in171;
input [7:0] in172;
input [7:0] in173;
input [7:0] in174;
input [7:0] in175;
input [7:0] in176;
input [7:0] in177;
input [7:0] in178;
input [7:0] in179;
input [7:0] in180;
input [7:0] in181;
input [7:0] in182;
input [7:0] in183;
input [7:0] in184;
input [7:0] in185;
input [7:0] in186;
input [7:0] in187;
input [7:0] in188;
input [7:0] in189;
input [7:0] in190;
input [7:0] in191;
input [7:0] in192;
input [7:0] in193;
input [7:0] in194;
input [7:0] in195;
input [7:0] in196;
input [7:0] in197;
input [7:0] in198;
input [7:0] in199;
input [7:0] in200;
input [7:0] in201;
input [7:0] in202;
input [7:0] in203;
input [7:0] in204;
input [7:0] in205;
input [7:0] in206;
input [7:0] in207;
input [7:0] in208;
input [7:0] in209;
input [7:0] in210;
input [7:0] in211;
input [7:0] in212;
input [7:0] in213;
input [7:0] in214;
input [7:0] in215;
input [7:0] in216;
input [7:0] in217;
input [7:0] in218;
input [7:0] in219;
input [7:0] in220;
input [7:0] in221;
input [7:0] in222;
input [7:0] in223;
input [7:0] in224;
input [7:0] in225;
input [7:0] in226;
input [7:0] in227;
input [7:0] in228;
input [7:0] in229;
input [7:0] in230;
input [7:0] in231;
input [7:0] in232;
input [7:0] in233;
input [7:0] in234;
input [7:0] in235;
input [7:0] in236;
input [7:0] in237;
input [7:0] in238;
input [7:0] in239;
input [7:0] in240;
input [7:0] in241;
input [7:0] in242;
input [7:0] in243;
input [7:0] in244;
input [7:0] in245;
input [7:0] in246;
input [7:0] in247;
input [7:0] in248;
input [7:0] in249;
input [7:0] in250;
input [7:0] in251;
input [7:0] in252;
input [7:0] in253;
input [7:0] in254;
input [7:0] in255;
input [7:0] in256;
input [7:0] in257;
input [7:0] in258;
input [7:0] in259;
input [7:0] in260;
input [7:0] in261;
input [7:0] in262;
input [7:0] in263;
input [7:0] in264;
input [7:0] in265;
input [7:0] in266;
input [7:0] in267;
input [7:0] in268;
input [7:0] in269;
input [7:0] in270;
input [7:0] in271;
input [7:0] in272;
input [7:0] in273;
input [7:0] in274;
input [7:0] in275;
input [7:0] in276;
input [7:0] in277;
input [7:0] in278;
input [7:0] in279;
input [7:0] in280;
input [7:0] in281;
input [7:0] in282;
input [7:0] in283;
input [7:0] in284;
input [7:0] in285;
input [7:0] in286;
input [7:0] in287;
input [7:0] in288;
input [7:0] in289;
input [7:0] in290;
input [7:0] in291;
input [7:0] in292;
input [7:0] in293;
input [7:0] in294;
input [7:0] in295;
input [7:0] in296;
input [7:0] in297;
input [7:0] in298;
input [7:0] in299;
input [7:0] in300;
input [7:0] in301;
input [7:0] in302;
input [7:0] in303;
input [7:0] in304;
input [7:0] in305;
input [7:0] in306;
input [7:0] in307;
input [7:0] in308;
input [7:0] in309;
input [7:0] in310;
input [7:0] in311;
input [7:0] in312;
input [7:0] in313;
input [7:0] in314;
input [7:0] in315;
input [7:0] in316;
input [7:0] in317;
input [7:0] in318;
input [7:0] in319;
input [7:0] in320;
input [7:0] in321;
input [7:0] in322;
input [7:0] in323;
input [7:0] in324;
input [7:0] in325;
input [7:0] in326;
input [7:0] in327;
input [7:0] in328;
input [7:0] in329;
input [7:0] in330;
input [7:0] in331;
input [7:0] in332;
input [7:0] in333;
input [7:0] in334;
input [7:0] in335;
input [7:0] in336;
input [7:0] in337;
input [7:0] in338;
input [7:0] in339;
input [7:0] in340;
input [7:0] in341;
input [7:0] in342;
input [7:0] in343;
input [7:0] in344;
input [7:0] in345;
input [7:0] in346;
input [7:0] in347;
input [7:0] in348;
input [7:0] in349;
input [7:0] in350;
input [7:0] in351;
input [7:0] in352;
input [7:0] in353;
input [7:0] in354;
input [7:0] in355;
input [7:0] in356;
input [7:0] in357;
input [7:0] in358;
input [7:0] in359;
input [7:0] in360;
input [7:0] in361;
input [7:0] in362;
input [7:0] in363;
input [7:0] in364;
input [7:0] in365;
input [7:0] in366;
input [7:0] in367;
input [7:0] in368;
input [7:0] in369;
input [7:0] in370;
input [7:0] in371;
input [7:0] in372;
input [7:0] in373;
input [7:0] in374;
input [7:0] in375;
input [7:0] in376;
input [7:0] in377;
input [7:0] in378;
input [7:0] in379;
input [7:0] in380;
input [7:0] in381;
input [7:0] in382;
input [7:0] in383;
input [7:0] in384;
input [7:0] in385;
input [7:0] in386;
input [7:0] in387;
input [7:0] in388;
input [7:0] in389;
input [7:0] in390;
input [7:0] in391;
input [7:0] in392;
input [7:0] in393;
input [7:0] in394;
input [7:0] in395;
input [7:0] in396;
input [7:0] in397;
input [7:0] in398;
input [7:0] in399;
input [7:0] in400;
input [7:0] in401;
input [7:0] in402;
input [7:0] in403;
input [7:0] in404;
input [7:0] in405;
input [7:0] in406;
input [7:0] in407;
input [7:0] in408;
input [7:0] in409;
input [7:0] in410;
input [7:0] in411;
input [7:0] in412;
input [7:0] in413;
input [7:0] in414;
input [7:0] in415;
input [7:0] in416;
input [7:0] in417;
input [7:0] in418;
input [7:0] in419;
input [7:0] in420;
input [7:0] in421;
input [7:0] in422;
input [7:0] in423;
input [7:0] in424;
input [7:0] in425;
input [7:0] in426;
input [7:0] in427;
input [7:0] in428;
input [7:0] in429;
input [7:0] in430;
input [7:0] in431;
input [7:0] in432;
input [7:0] in433;
input [7:0] in434;
input [7:0] in435;
input [7:0] in436;
input [7:0] in437;
input [7:0] in438;
input [7:0] in439;
input [7:0] in440;
input [7:0] in441;
input [7:0] in442;
input [7:0] in443;
input [7:0] in444;
input [7:0] in445;
input [7:0] in446;
input [7:0] in447;
input [7:0] in448;
input [7:0] in449;
input [7:0] in450;
input [7:0] in451;
input [7:0] in452;
input [7:0] in453;
input [7:0] in454;
input [7:0] in455;
input [7:0] in456;
input [7:0] in457;
input [7:0] in458;
input [7:0] in459;
input [7:0] in460;
input [7:0] in461;
input [7:0] in462;
input [7:0] in463;
input [7:0] in464;
input [7:0] in465;
input [7:0] in466;
input [7:0] in467;
input [7:0] in468;
input [7:0] in469;
input [7:0] in470;
input [7:0] in471;
input [7:0] in472;
input [7:0] in473;
input [7:0] in474;
input [7:0] in475;
input [7:0] in476;
input [7:0] in477;
input [7:0] in478;
input [7:0] in479;
input [7:0] in480;
input [7:0] in481;
input [7:0] in482;
input [7:0] in483;
input [7:0] in484;
input [7:0] in485;
input [7:0] in486;
input [7:0] in487;
input [7:0] in488;
input [7:0] in489;
input [7:0] in490;
input [7:0] in491;
input [7:0] in492;
input [7:0] in493;
input [7:0] in494;
input [7:0] in495;
input [7:0] in496;
input [7:0] in497;
input [7:0] in498;
input [7:0] in499;
input [7:0] in500;
input [7:0] in501;
input [7:0] in502;
input [7:0] in503;
input [7:0] in504;
input [7:0] in505;
input [7:0] in506;
input [7:0] in507;
input [7:0] in508;
input [7:0] in509;
input [7:0] in510;
input [7:0] in511;
input [7:0] in512;
input [7:0] in513;
input [7:0] in514;
input [7:0] in515;
input [7:0] in516;
input [7:0] in517;
input [7:0] in518;
input [7:0] in519;
input [7:0] in520;
input [7:0] in521;
input [7:0] in522;
input [7:0] in523;
input [7:0] in524;
input [7:0] in525;
input [7:0] in526;
input [7:0] in527;
input [7:0] in528;
input [7:0] in529;
input [7:0] in530;
input [7:0] in531;
input [7:0] in532;
input [7:0] in533;
input [7:0] in534;
input [7:0] in535;
input [7:0] in536;
input [7:0] in537;
input [7:0] in538;
input [7:0] in539;
input [7:0] in540;
input [7:0] in541;
input [7:0] in542;
input [7:0] in543;
input [7:0] in544;
input [7:0] in545;
input [7:0] in546;
input [7:0] in547;
input [7:0] in548;
input [7:0] in549;
input [7:0] in550;
input [7:0] in551;
input [7:0] in552;
input [7:0] in553;
input [7:0] in554;
input [7:0] in555;
input [7:0] in556;
input [7:0] in557;
input [7:0] in558;
input [7:0] in559;
input [7:0] in560;
input [7:0] in561;
input [7:0] in562;
input [7:0] in563;
input [7:0] in564;
input [7:0] in565;
input [7:0] in566;
input [7:0] in567;
input [7:0] in568;
input [7:0] in569;
input [7:0] in570;
input [7:0] in571;
input [7:0] in572;
input [7:0] in573;
input [7:0] in574;
input [7:0] in575;
input [7:0] in576;
input [7:0] in577;
input [7:0] in578;
input [7:0] in579;
input [7:0] in580;
input [7:0] in581;
input [7:0] in582;
input [7:0] in583;
input [7:0] in584;
input [7:0] in585;
input [7:0] in586;
input [7:0] in587;
input [7:0] in588;
input [7:0] in589;
input [7:0] in590;
input [7:0] in591;
input [7:0] in592;
input [7:0] in593;
input [7:0] in594;
input [7:0] in595;
input [7:0] in596;
input [7:0] in597;
input [7:0] in598;
input [7:0] in599;
input [7:0] in600;
input [7:0] in601;
input [7:0] in602;
input [7:0] in603;
input [7:0] in604;
input [7:0] in605;
input [7:0] in606;
input [7:0] in607;
input [7:0] in608;
input [7:0] in609;
input [7:0] in610;
input [7:0] in611;
input [7:0] in612;
input [7:0] in613;
input [7:0] in614;
input [7:0] in615;
input [7:0] in616;
input [7:0] in617;
input [7:0] in618;
input [7:0] in619;
input [7:0] in620;
input [7:0] in621;
input [7:0] in622;
input [7:0] in623;
input [7:0] in624;
input [7:0] in625;
input [7:0] in626;
input [7:0] in627;
input [7:0] in628;
input [7:0] in629;
input [7:0] in630;
input [7:0] in631;
input [7:0] in632;
input [7:0] in633;
input [7:0] in634;
input [7:0] in635;
input [7:0] in636;
input [7:0] in637;
input [7:0] in638;
input [7:0] in639;
input [7:0] in640;
input [7:0] in641;
input [7:0] in642;
input [7:0] in643;
input [7:0] in644;
input [7:0] in645;
input [7:0] in646;
input [7:0] in647;
input [7:0] in648;
input [7:0] in649;
input [7:0] in650;
input [7:0] in651;
input [7:0] in652;
input [7:0] in653;
input [7:0] in654;
input [7:0] in655;
input [7:0] in656;
input [7:0] in657;
input [7:0] in658;
input [7:0] in659;
input [7:0] in660;
input [7:0] in661;
input [7:0] in662;
input [7:0] in663;
input [7:0] in664;
input [7:0] in665;
input [7:0] in666;
input [7:0] in667;
input [7:0] in668;
input [7:0] in669;
input [7:0] in670;
input [7:0] in671;
input [7:0] in672;
input [7:0] in673;
input [7:0] in674;
input [7:0] in675;
input [7:0] in676;
input [7:0] in677;
input [7:0] in678;
input [7:0] in679;
input [7:0] in680;
input [7:0] in681;
input [7:0] in682;
input [7:0] in683;
input [7:0] in684;
input [7:0] in685;
input [7:0] in686;
input [7:0] in687;
input [7:0] in688;
input [7:0] in689;
input [7:0] in690;
input [7:0] in691;
input [7:0] in692;
input [7:0] in693;
input [7:0] in694;
input [7:0] in695;
input [7:0] in696;
input [7:0] in697;
input [7:0] in698;
input [7:0] in699;
input [7:0] in700;
input [7:0] in701;
input [7:0] in702;
input [7:0] in703;
input [7:0] in704;
input [7:0] in705;
input [7:0] in706;
input [7:0] in707;
input [7:0] in708;
input [7:0] in709;
input [7:0] in710;
input [7:0] in711;
input [7:0] in712;
input [7:0] in713;
input [7:0] in714;
input [7:0] in715;
input [7:0] in716;
input [7:0] in717;
input [7:0] in718;
input [7:0] in719;
input [7:0] in720;
input [7:0] in721;
input [7:0] in722;
input [7:0] in723;
input [7:0] in724;
input [7:0] in725;
input [7:0] in726;
input [7:0] in727;
input [7:0] in728;
input [7:0] in729;
input [7:0] in730;
input [7:0] in731;
input [7:0] in732;
input [7:0] in733;
input [7:0] in734;
input [7:0] in735;
input [7:0] in736;
input [7:0] in737;
input [7:0] in738;
input [7:0] in739;
input [7:0] in740;
input [7:0] in741;
input [7:0] in742;
input [7:0] in743;
input [7:0] in744;
input [7:0] in745;
input [7:0] in746;
input [7:0] in747;
input [7:0] in748;
input [7:0] in749;
input [7:0] in750;
input [7:0] in751;
input [7:0] in752;
input [7:0] in753;
input [7:0] in754;
input [7:0] in755;
input [7:0] in756;
input [7:0] in757;
input [7:0] in758;
input [7:0] in759;
input [7:0] in760;
input [7:0] in761;
input [7:0] in762;
input [7:0] in763;
input [7:0] in764;
input [7:0] in765;
input [7:0] in766;
input [7:0] in767;
input [7:0] in768;
input [7:0] in769;
input [7:0] in770;
input [7:0] in771;
input [7:0] in772;
input [7:0] in773;
input [7:0] in774;
input [7:0] in775;
input [7:0] in776;
input [7:0] in777;
input [7:0] in778;
input [7:0] in779;
input [7:0] in780;
input [7:0] in781;
input [7:0] in782;
input [7:0] in783;

input [7:0] weight0;
input [7:0] weight1;
input [7:0] weight2;
input [7:0] weight3;
input [7:0] weight4;
input [7:0] weight5;
input [7:0] weight6;
input [7:0] weight7;
input [7:0] weight8;
input [7:0] weight9;
input [7:0] weight10;
input [7:0] weight11;
input [7:0] weight12;
input [7:0] weight13;
input [7:0] weight14;
input [7:0] weight15;
input [7:0] weight16;
input [7:0] weight17;
input [7:0] weight18;
input [7:0] weight19;
input [7:0] weight20;
input [7:0] weight21;
input [7:0] weight22;
input [7:0] weight23;
input [7:0] weight24;

input [7:0] bias;
input clk;


 output [7:0] conv0;
output [7:0] conv1;
output [7:0] conv2;
output [7:0] conv3;
output [7:0] conv4;
output [7:0] conv5;
output [7:0] conv6;
output [7:0] conv7;
output [7:0] conv8;
output [7:0] conv9;
output [7:0] conv10;
output [7:0] conv11;
output [7:0] conv12;
output [7:0] conv13;
output [7:0] conv14;
output [7:0] conv15;
output [7:0] conv16;
output [7:0] conv17;
output [7:0] conv18;
output [7:0] conv19;
output [7:0] conv20;
output [7:0] conv21;
output [7:0] conv22;
output [7:0] conv23;
output [7:0] conv24;
output [7:0] conv25;
output [7:0] conv26;
output [7:0] conv27;
output [7:0] conv28;
output [7:0] conv29;
output [7:0] conv30;
output [7:0] conv31;
output [7:0] conv32;
output [7:0] conv33;
output [7:0] conv34;
output [7:0] conv35;
output [7:0] conv36;
output [7:0] conv37;
output [7:0] conv38;
output [7:0] conv39;
output [7:0] conv40;
output [7:0] conv41;
output [7:0] conv42;
output [7:0] conv43;
output [7:0] conv44;
output [7:0] conv45;
output [7:0] conv46;
output [7:0] conv47;
output [7:0] conv48;
output [7:0] conv49;
output [7:0] conv50;
output [7:0] conv51;
output [7:0] conv52;
output [7:0] conv53;
output [7:0] conv54;
output [7:0] conv55;
output [7:0] conv56;
output [7:0] conv57;
output [7:0] conv58;
output [7:0] conv59;
output [7:0] conv60;
output [7:0] conv61;
output [7:0] conv62;
output [7:0] conv63;
output [7:0] conv64;
output [7:0] conv65;
output [7:0] conv66;
output [7:0] conv67;
output [7:0] conv68;
output [7:0] conv69;
output [7:0] conv70;
output [7:0] conv71;
output [7:0] conv72;
output [7:0] conv73;
output [7:0] conv74;
output [7:0] conv75;
output [7:0] conv76;
output [7:0] conv77;
output [7:0] conv78;
output [7:0] conv79;
output [7:0] conv80;
output [7:0] conv81;
output [7:0] conv82;
output [7:0] conv83;
output [7:0] conv84;
output [7:0] conv85;
output [7:0] conv86;
output [7:0] conv87;
output [7:0] conv88;
output [7:0] conv89;
output [7:0] conv90;
output [7:0] conv91;
output [7:0] conv92;
output [7:0] conv93;
output [7:0] conv94;
output [7:0] conv95;
output [7:0] conv96;
output [7:0] conv97;
output [7:0] conv98;
output [7:0] conv99;
output [7:0] conv100;
output [7:0] conv101;
output [7:0] conv102;
output [7:0] conv103;
output [7:0] conv104;
output [7:0] conv105;
output [7:0] conv106;
output [7:0] conv107;
output [7:0] conv108;
output [7:0] conv109;
output [7:0] conv110;
output [7:0] conv111;
output [7:0] conv112;
output [7:0] conv113;
output [7:0] conv114;
output [7:0] conv115;
output [7:0] conv116;
output [7:0] conv117;
output [7:0] conv118;
output [7:0] conv119;
output [7:0] conv120;
output [7:0] conv121;
output [7:0] conv122;
output [7:0] conv123;
output [7:0] conv124;
output [7:0] conv125;
output [7:0] conv126;
output [7:0] conv127;
output [7:0] conv128;
output [7:0] conv129;
output [7:0] conv130;
output [7:0] conv131;
output [7:0] conv132;
output [7:0] conv133;
output [7:0] conv134;
output [7:0] conv135;
output [7:0] conv136;
output [7:0] conv137;
output [7:0] conv138;
output [7:0] conv139;
output [7:0] conv140;
output [7:0] conv141;
output [7:0] conv142;
output [7:0] conv143;
output [7:0] conv144;
output [7:0] conv145;
output [7:0] conv146;
output [7:0] conv147;
output [7:0] conv148;
output [7:0] conv149;
output [7:0] conv150;
output [7:0] conv151;
output [7:0] conv152;
output [7:0] conv153;
output [7:0] conv154;
output [7:0] conv155;
output [7:0] conv156;
output [7:0] conv157;
output [7:0] conv158;
output [7:0] conv159;
output [7:0] conv160;
output [7:0] conv161;
output [7:0] conv162;
output [7:0] conv163;
output [7:0] conv164;
output [7:0] conv165;
output [7:0] conv166;
output [7:0] conv167;
output [7:0] conv168;
output [7:0] conv169;
output [7:0] conv170;
output [7:0] conv171;
output [7:0] conv172;
output [7:0] conv173;
output [7:0] conv174;
output [7:0] conv175;
output [7:0] conv176;
output [7:0] conv177;
output [7:0] conv178;
output [7:0] conv179;
output [7:0] conv180;
output [7:0] conv181;
output [7:0] conv182;
output [7:0] conv183;
output [7:0] conv184;
output [7:0] conv185;
output [7:0] conv186;
output [7:0] conv187;
output [7:0] conv188;
output [7:0] conv189;
output [7:0] conv190;
output [7:0] conv191;
output [7:0] conv192;
output [7:0] conv193;
output [7:0] conv194;
output [7:0] conv195;
output [7:0] conv196;
output [7:0] conv197;
output [7:0] conv198;
output [7:0] conv199;
output [7:0] conv200;
output [7:0] conv201;
output [7:0] conv202;
output [7:0] conv203;
output [7:0] conv204;
output [7:0] conv205;
output [7:0] conv206;
output [7:0] conv207;
output [7:0] conv208;
output [7:0] conv209;
output [7:0] conv210;
output [7:0] conv211;
output [7:0] conv212;
output [7:0] conv213;
output [7:0] conv214;
output [7:0] conv215;
output [7:0] conv216;
output [7:0] conv217;
output [7:0] conv218;
output [7:0] conv219;
output [7:0] conv220;
output [7:0] conv221;
output [7:0] conv222;
output [7:0] conv223;
output [7:0] conv224;
output [7:0] conv225;
output [7:0] conv226;
output [7:0] conv227;
output [7:0] conv228;
output [7:0] conv229;
output [7:0] conv230;
output [7:0] conv231;
output [7:0] conv232;
output [7:0] conv233;
output [7:0] conv234;
output [7:0] conv235;
output [7:0] conv236;
output [7:0] conv237;
output [7:0] conv238;
output [7:0] conv239;
output [7:0] conv240;
output [7:0] conv241;
output [7:0] conv242;
output [7:0] conv243;
output [7:0] conv244;
output [7:0] conv245;
output [7:0] conv246;
output [7:0] conv247;
output [7:0] conv248;
output [7:0] conv249;
output [7:0] conv250;
output [7:0] conv251;
output [7:0] conv252;
output [7:0] conv253;
output [7:0] conv254;
output [7:0] conv255;
output [7:0] conv256;
output [7:0] conv257;
output [7:0] conv258;
output [7:0] conv259;
output [7:0] conv260;
output [7:0] conv261;
output [7:0] conv262;
output [7:0] conv263;
output [7:0] conv264;
output [7:0] conv265;
output [7:0] conv266;
output [7:0] conv267;
output [7:0] conv268;
output [7:0] conv269;
output [7:0] conv270;
output [7:0] conv271;
output [7:0] conv272;
output [7:0] conv273;
output [7:0] conv274;
output [7:0] conv275;
output [7:0] conv276;
output [7:0] conv277;
output [7:0] conv278;
output [7:0] conv279;
output [7:0] conv280;
output [7:0] conv281;
output [7:0] conv282;
output [7:0] conv283;
output [7:0] conv284;
output [7:0] conv285;
output [7:0] conv286;
output [7:0] conv287;
output [7:0] conv288;
output [7:0] conv289;
output [7:0] conv290;
output [7:0] conv291;
output [7:0] conv292;
output [7:0] conv293;
output [7:0] conv294;
output [7:0] conv295;
output [7:0] conv296;
output [7:0] conv297;
output [7:0] conv298;
output [7:0] conv299;
output [7:0] conv300;
output [7:0] conv301;
output [7:0] conv302;
output [7:0] conv303;
output [7:0] conv304;
output [7:0] conv305;
output [7:0] conv306;
output [7:0] conv307;
output [7:0] conv308;
output [7:0] conv309;
output [7:0] conv310;
output [7:0] conv311;
output [7:0] conv312;
output [7:0] conv313;
output [7:0] conv314;
output [7:0] conv315;
output [7:0] conv316;
output [7:0] conv317;
output [7:0] conv318;
output [7:0] conv319;
output [7:0] conv320;
output [7:0] conv321;
output [7:0] conv322;
output [7:0] conv323;
output [7:0] conv324;
output [7:0] conv325;
output [7:0] conv326;
output [7:0] conv327;
output [7:0] conv328;
output [7:0] conv329;
output [7:0] conv330;
output [7:0] conv331;
output [7:0] conv332;
output [7:0] conv333;
output [7:0] conv334;
output [7:0] conv335;
output [7:0] conv336;
output [7:0] conv337;
output [7:0] conv338;
output [7:0] conv339;
output [7:0] conv340;
output [7:0] conv341;
output [7:0] conv342;
output [7:0] conv343;
output [7:0] conv344;
output [7:0] conv345;
output [7:0] conv346;
output [7:0] conv347;
output [7:0] conv348;
output [7:0] conv349;
output [7:0] conv350;
output [7:0] conv351;
output [7:0] conv352;
output [7:0] conv353;
output [7:0] conv354;
output [7:0] conv355;
output [7:0] conv356;
output [7:0] conv357;
output [7:0] conv358;
output [7:0] conv359;
output [7:0] conv360;
output [7:0] conv361;
output [7:0] conv362;
output [7:0] conv363;
output [7:0] conv364;
output [7:0] conv365;
output [7:0] conv366;
output [7:0] conv367;
output [7:0] conv368;
output [7:0] conv369;
output [7:0] conv370;
output [7:0] conv371;
output [7:0] conv372;
output [7:0] conv373;
output [7:0] conv374;
output [7:0] conv375;
output [7:0] conv376;
output [7:0] conv377;
output [7:0] conv378;
output [7:0] conv379;
output [7:0] conv380;
output [7:0] conv381;
output [7:0] conv382;
output [7:0] conv383;
output [7:0] conv384;
output [7:0] conv385;
output [7:0] conv386;
output [7:0] conv387;
output [7:0] conv388;
output [7:0] conv389;
output [7:0] conv390;
output [7:0] conv391;
output [7:0] conv392;
output [7:0] conv393;
output [7:0] conv394;
output [7:0] conv395;
output [7:0] conv396;
output [7:0] conv397;
output [7:0] conv398;
output [7:0] conv399;
output [7:0] conv400;
output [7:0] conv401;
output [7:0] conv402;
output [7:0] conv403;
output [7:0] conv404;
output [7:0] conv405;
output [7:0] conv406;
output [7:0] conv407;
output [7:0] conv408;
output [7:0] conv409;
output [7:0] conv410;
output [7:0] conv411;
output [7:0] conv412;
output [7:0] conv413;
output [7:0] conv414;
output [7:0] conv415;
output [7:0] conv416;
output [7:0] conv417;
output [7:0] conv418;
output [7:0] conv419;
output [7:0] conv420;
output [7:0] conv421;
output [7:0] conv422;
output [7:0] conv423;
output [7:0] conv424;
output [7:0] conv425;
output [7:0] conv426;
output [7:0] conv427;
output [7:0] conv428;
output [7:0] conv429;
output [7:0] conv430;
output [7:0] conv431;
output [7:0] conv432;
output [7:0] conv433;
output [7:0] conv434;
output [7:0] conv435;
output [7:0] conv436;
output [7:0] conv437;
output [7:0] conv438;
output [7:0] conv439;
output [7:0] conv440;
output [7:0] conv441;
output [7:0] conv442;
output [7:0] conv443;
output [7:0] conv444;
output [7:0] conv445;
output [7:0] conv446;
output [7:0] conv447;
output [7:0] conv448;
output [7:0] conv449;
output [7:0] conv450;
output [7:0] conv451;
output [7:0] conv452;
output [7:0] conv453;
output [7:0] conv454;
output [7:0] conv455;
output [7:0] conv456;
output [7:0] conv457;
output [7:0] conv458;
output [7:0] conv459;
output [7:0] conv460;
output [7:0] conv461;
output [7:0] conv462;
output [7:0] conv463;
output [7:0] conv464;
output [7:0] conv465;
output [7:0] conv466;
output [7:0] conv467;
output [7:0] conv468;
output [7:0] conv469;
output [7:0] conv470;
output [7:0] conv471;
output [7:0] conv472;
output [7:0] conv473;
output [7:0] conv474;
output [7:0] conv475;
output [7:0] conv476;
output [7:0] conv477;
output [7:0] conv478;
output [7:0] conv479;
output [7:0] conv480;
output [7:0] conv481;
output [7:0] conv482;
output [7:0] conv483;
output [7:0] conv484;
output [7:0] conv485;
output [7:0] conv486;
output [7:0] conv487;
output [7:0] conv488;
output [7:0] conv489;
output [7:0] conv490;
output [7:0] conv491;
output [7:0] conv492;
output [7:0] conv493;
output [7:0] conv494;
output [7:0] conv495;
output [7:0] conv496;
output [7:0] conv497;
output [7:0] conv498;
output [7:0] conv499;
output [7:0] conv500;
output [7:0] conv501;
output [7:0] conv502;
output [7:0] conv503;
output [7:0] conv504;
output [7:0] conv505;
output [7:0] conv506;
output [7:0] conv507;
output [7:0] conv508;
output [7:0] conv509;
output [7:0] conv510;
output [7:0] conv511;
output [7:0] conv512;
output [7:0] conv513;
output [7:0] conv514;
output [7:0] conv515;
output [7:0] conv516;
output [7:0] conv517;
output [7:0] conv518;
output [7:0] conv519;
output [7:0] conv520;
output [7:0] conv521;
output [7:0] conv522;
output [7:0] conv523;
output [7:0] conv524;
output [7:0] conv525;
output [7:0] conv526;
output [7:0] conv527;
output [7:0] conv528;
output [7:0] conv529;
output [7:0] conv530;
output [7:0] conv531;
output [7:0] conv532;
output [7:0] conv533;
output [7:0] conv534;
output [7:0] conv535;
output [7:0] conv536;
output [7:0] conv537;
output [7:0] conv538;
output [7:0] conv539;
output [7:0] conv540;
output [7:0] conv541;
output [7:0] conv542;
output [7:0] conv543;
output [7:0] conv544;
output [7:0] conv545;
output [7:0] conv546;
output [7:0] conv547;
output [7:0] conv548;
output [7:0] conv549;
output [7:0] conv550;
output [7:0] conv551;
output [7:0] conv552;
output [7:0] conv553;
output [7:0] conv554;
output [7:0] conv555;
output [7:0] conv556;
output [7:0] conv557;
output [7:0] conv558;
output [7:0] conv559;
output [7:0] conv560;
output [7:0] conv561;
output [7:0] conv562;
output [7:0] conv563;
output [7:0] conv564;
output [7:0] conv565;
output [7:0] conv566;
output [7:0] conv567;
output [7:0] conv568;
output [7:0] conv569;
output [7:0] conv570;
output [7:0] conv571;
output [7:0] conv572;
output [7:0] conv573;
output [7:0] conv574;
output [7:0] conv575;

wire [7:0] mux0;
wire [7:0] mux1;
wire [7:0] mux2;
wire [7:0] mux3;
wire [7:0] mux4;
wire [7:0] mux5;
wire [7:0] mux6;
wire [7:0] mux7;
wire [7:0] mux8;
wire [7:0] mux9;
wire [7:0] mux10;
wire [7:0] mux11;
wire [7:0] mux12;
wire [7:0] mux13;
wire [7:0] mux14;
wire [7:0] mux15;
wire [7:0] mux16;
wire [7:0] mux17;
wire [7:0] mux18;
wire [7:0] mux19;
wire [7:0] mux20;
wire [7:0] mux21;
wire [7:0] mux22;
wire [7:0] mux23;
wire [7:0] mux24;
wire [7:0] mux25;
wire [7:0] mux26;
wire [7:0] mux27;
wire [7:0] mux28;
wire [7:0] mux29;
wire [7:0] mux30;
wire [7:0] mux31;
wire [7:0] mux32;
wire [7:0] mux33;
wire [7:0] mux34;
wire [7:0] mux35;
wire [7:0] mux36;
wire [7:0] mux37;
wire [7:0] mux38;
wire [7:0] mux39;
wire [7:0] mux40;
wire [7:0] mux41;
wire [7:0] mux42;
wire [7:0] mux43;
wire [7:0] mux44;
wire [7:0] mux45;
wire [7:0] mux46;
wire [7:0] mux47;
wire [7:0] mux48;
wire [7:0] mux49;
wire [7:0] mux50;
wire [7:0] mux51;
wire [7:0] mux52;
wire [7:0] mux53;
wire [7:0] mux54;
wire [7:0] mux55;
wire [7:0] mux56;
wire [7:0] mux57;
wire [7:0] mux58;
wire [7:0] mux59;
wire [7:0] mux60;
wire [7:0] mux61;
wire [7:0] mux62;
wire [7:0] mux63;
wire [7:0] mux64;
wire [7:0] mux65;
wire [7:0] mux66;
wire [7:0] mux67;
wire [7:0] mux68;
wire [7:0] mux69;
wire [7:0] mux70;
wire [7:0] mux71;
wire [7:0] mux72;
wire [7:0] mux73;
wire [7:0] mux74;
wire [7:0] mux75;
wire [7:0] mux76;
wire [7:0] mux77;
wire [7:0] mux78;
wire [7:0] mux79;
wire [7:0] mux80;
wire [7:0] mux81;
wire [7:0] mux82;
wire [7:0] mux83;
wire [7:0] mux84;
wire [7:0] mux85;
wire [7:0] mux86;
wire [7:0] mux87;
wire [7:0] mux88;
wire [7:0] mux89;
wire [7:0] mux90;
wire [7:0] mux91;
wire [7:0] mux92;
wire [7:0] mux93;
wire [7:0] mux94;
wire [7:0] mux95;
wire [7:0] mux96;
wire [7:0] mux97;
wire [7:0] mux98;
wire [7:0] mux99;
wire [7:0] mux100;
wire [7:0] mux101;
wire [7:0] mux102;
wire [7:0] mux103;
wire [7:0] mux104;
wire [7:0] mux105;
wire [7:0] mux106;
wire [7:0] mux107;
wire [7:0] mux108;
wire [7:0] mux109;
wire [7:0] mux110;
wire [7:0] mux111;
wire [7:0] mux112;
wire [7:0] mux113;
wire [7:0] mux114;
wire [7:0] mux115;
wire [7:0] mux116;
wire [7:0] mux117;
wire [7:0] mux118;
wire [7:0] mux119;
wire [7:0] mux120;
wire [7:0] mux121;
wire [7:0] mux122;
wire [7:0] mux123;
wire [7:0] mux124;
wire [7:0] mux125;
wire [7:0] mux126;
wire [7:0] mux127;
wire [7:0] mux128;
wire [7:0] mux129;
wire [7:0] mux130;
wire [7:0] mux131;
wire [7:0] mux132;
wire [7:0] mux133;
wire [7:0] mux134;
wire [7:0] mux135;
wire [7:0] mux136;
wire [7:0] mux137;
wire [7:0] mux138;
wire [7:0] mux139;
wire [7:0] mux140;
wire [7:0] mux141;
wire [7:0] mux142;
wire [7:0] mux143;
wire [7:0] mux144;
wire [7:0] mux145;
wire [7:0] mux146;
wire [7:0] mux147;
wire [7:0] mux148;
wire [7:0] mux149;
wire [7:0] mux150;
wire [7:0] mux151;
wire [7:0] mux152;
wire [7:0] mux153;
wire [7:0] mux154;
wire [7:0] mux155;
wire [7:0] mux156;
wire [7:0] mux157;
wire [7:0] mux158;
wire [7:0] mux159;
wire [7:0] mux160;
wire [7:0] mux161;
wire [7:0] mux162;
wire [7:0] mux163;
wire [7:0] mux164;
wire [7:0] mux165;
wire [7:0] mux166;
wire [7:0] mux167;
wire [7:0] mux168;
wire [7:0] mux169;
wire [7:0] mux170;
wire [7:0] mux171;
wire [7:0] mux172;
wire [7:0] mux173;
wire [7:0] mux174;
wire [7:0] mux175;
wire [7:0] mux176;
wire [7:0] mux177;
wire [7:0] mux178;
wire [7:0] mux179;
wire [7:0] mux180;
wire [7:0] mux181;
wire [7:0] mux182;
wire [7:0] mux183;
wire [7:0] mux184;
wire [7:0] mux185;
wire [7:0] mux186;
wire [7:0] mux187;
wire [7:0] mux188;
wire [7:0] mux189;
wire [7:0] mux190;
wire [7:0] mux191;
wire [7:0] mux192;
wire [7:0] mux193;
wire [7:0] mux194;
wire [7:0] mux195;
wire [7:0] mux196;
wire [7:0] mux197;
wire [7:0] mux198;
wire [7:0] mux199;
wire [7:0] mux200;
wire [7:0] mux201;
wire [7:0] mux202;
wire [7:0] mux203;
wire [7:0] mux204;
wire [7:0] mux205;
wire [7:0] mux206;
wire [7:0] mux207;
wire [7:0] mux208;
wire [7:0] mux209;
wire [7:0] mux210;
wire [7:0] mux211;
wire [7:0] mux212;
wire [7:0] mux213;
wire [7:0] mux214;
wire [7:0] mux215;
wire [7:0] mux216;
wire [7:0] mux217;
wire [7:0] mux218;
wire [7:0] mux219;
wire [7:0] mux220;
wire [7:0] mux221;
wire [7:0] mux222;
wire [7:0] mux223;
wire [7:0] mux224;
wire [7:0] mux225;
wire [7:0] mux226;
wire [7:0] mux227;
wire [7:0] mux228;
wire [7:0] mux229;
wire [7:0] mux230;
wire [7:0] mux231;
wire [7:0] mux232;
wire [7:0] mux233;
wire [7:0] mux234;
wire [7:0] mux235;
wire [7:0] mux236;
wire [7:0] mux237;
wire [7:0] mux238;
wire [7:0] mux239;
wire [7:0] mux240;
wire [7:0] mux241;
wire [7:0] mux242;
wire [7:0] mux243;
wire [7:0] mux244;
wire [7:0] mux245;
wire [7:0] mux246;
wire [7:0] mux247;
wire [7:0] mux248;
wire [7:0] mux249;
wire [7:0] mux250;
wire [7:0] mux251;
wire [7:0] mux252;
wire [7:0] mux253;
wire [7:0] mux254;
wire [7:0] mux255;
wire [7:0] mux256;
wire [7:0] mux257;
wire [7:0] mux258;
wire [7:0] mux259;
wire [7:0] mux260;
wire [7:0] mux261;
wire [7:0] mux262;
wire [7:0] mux263;
wire [7:0] mux264;
wire [7:0] mux265;
wire [7:0] mux266;
wire [7:0] mux267;
wire [7:0] mux268;
wire [7:0] mux269;
wire [7:0] mux270;
wire [7:0] mux271;
wire [7:0] mux272;
wire [7:0] mux273;
wire [7:0] mux274;
wire [7:0] mux275;
wire [7:0] mux276;
wire [7:0] mux277;
wire [7:0] mux278;
wire [7:0] mux279;


 wire [7:0] muxin0;
wire [7:0] muxin1;
wire [7:0] muxin2;
wire [7:0] muxin3;
wire [7:0] muxin4;
wire [7:0] muxin5;
wire [7:0] muxin6;
wire [7:0] muxin7;
wire [7:0] muxin8;
wire [7:0] muxin9;
wire [7:0] muxin10;
wire [7:0] muxin11;
wire [7:0] muxin12;
wire [7:0] muxin13;
wire [7:0] muxin14;
wire [7:0] muxin15;
wire [7:0] muxin16;
wire [7:0] muxin17;
wire [7:0] muxin18;
wire [7:0] muxin19;
wire [7:0] muxin20;
wire [7:0] muxin21;
wire [7:0] muxin22;
wire [7:0] muxin23;
wire [7:0] muxin24;
wire [7:0] muxin25;
wire [7:0] muxin26;
wire [7:0] muxin27;
wire [7:0] muxin28;
wire [7:0] muxin29;
wire [7:0] muxin30;
wire [7:0] muxin31;
wire [7:0] muxin32;
wire [7:0] muxin33;
wire [7:0] muxin34;
wire [7:0] muxin35;
wire [7:0] muxin36;
wire [7:0] muxin37;
wire [7:0] muxin38;
wire [7:0] muxin39;
wire [7:0] muxin40;
wire [7:0] muxin41;
wire [7:0] muxin42;
wire [7:0] muxin43;
wire [7:0] muxin44;
wire [7:0] muxin45;
wire [7:0] muxin46;
wire [7:0] muxin47;
wire [7:0] muxin48;
wire [7:0] muxin49;
wire [7:0] muxin50;
wire [7:0] muxin51;
wire [7:0] muxin52;
wire [7:0] muxin53;
wire [7:0] muxin54;
wire [7:0] muxin55;
wire [7:0] muxin56;
wire [7:0] muxin57;
wire [7:0] muxin58;
wire [7:0] muxin59;
wire [7:0] muxin60;
wire [7:0] muxin61;
wire [7:0] muxin62;
wire [7:0] muxin63;
wire [7:0] muxin64;
wire [7:0] muxin65;
wire [7:0] muxin66;
wire [7:0] muxin67;
wire [7:0] muxin68;
wire [7:0] muxin69;
wire [7:0] muxin70;
wire [7:0] muxin71;
wire [7:0] muxin72;
wire [7:0] muxin73;
wire [7:0] muxin74;
wire [7:0] muxin75;
wire [7:0] muxin76;
wire [7:0] muxin77;
wire [7:0] muxin78;
wire [7:0] muxin79;
wire [7:0] muxin80;
wire [7:0] muxin81;
wire [7:0] muxin82;
wire [7:0] muxin83;
wire [7:0] muxin84;
wire [7:0] muxin85;
wire [7:0] muxin86;
wire [7:0] muxin87;
wire [7:0] muxin88;
wire [7:0] muxin89;
wire [7:0] muxin90;
wire [7:0] muxin91;
wire [7:0] muxin92;
wire [7:0] muxin93;
wire [7:0] muxin94;
wire [7:0] muxin95;
wire [7:0] muxin96;
wire [7:0] muxin97;
wire [7:0] muxin98;
wire [7:0] muxin99;
wire [7:0] muxin100;
wire [7:0] muxin101;
wire [7:0] muxin102;
wire [7:0] muxin103;
wire [7:0] muxin104;
wire [7:0] muxin105;
wire [7:0] muxin106;
wire [7:0] muxin107;
wire [7:0] muxin108;
wire [7:0] muxin109;
wire [7:0] muxin110;
wire [7:0] muxin111;
wire [7:0] muxin112;
wire [7:0] muxin113;
wire [7:0] muxin114;
wire [7:0] muxin115;
wire [7:0] muxin116;
wire [7:0] muxin117;
wire [7:0] muxin118;
wire [7:0] muxin119;
wire [7:0] muxin120;
wire [7:0] muxin121;
wire [7:0] muxin122;
wire [7:0] muxin123;
wire [7:0] muxin124;
wire [7:0] muxin125;
wire [7:0] muxin126;
wire [7:0] muxin127;
wire [7:0] muxin128;
wire [7:0] muxin129;
wire [7:0] muxin130;
wire [7:0] muxin131;
wire [7:0] muxin132;
wire [7:0] muxin133;
wire [7:0] muxin134;
wire [7:0] muxin135;
wire [7:0] muxin136;
wire [7:0] muxin137;
wire [7:0] muxin138;
wire [7:0] muxin139;
wire [7:0] muxin140;
wire [7:0] muxin141;
wire [7:0] muxin142;
wire [7:0] muxin143;

reg [1:0] sel;
reg [2:0] state;
reg [2:0] next_state;


always @(posedge start or posedge clk)
begin
	//$monitor(ready);
	if (start) begin
		next_state <= 3'b111;
		ready <= 0;
	end
	else
	begin
	state <= next_state;
	end
	case ({state})
		{3'b111}:
			begin
				sel <= 2'b00;
				next_state <= 3'b001;
			end
		{3'b001}:
			begin
				sel <= 2'b00;
				next_state <= 3'b010;
			end
		{3'b010}:
			begin
				sel <= 2'b01;
				next_state <= 3'b011;
			end
		{3'b011}:
			begin
				sel <= 2'b10;
				next_state <= 3'b100;
			end
		{3'b100}:
			begin
				sel <= 2'b11;
				next_state <= 3'b101;
				ready <= 0;
			end
		{3'b101}:
			begin
				sel <= 2'b00;
				next_state <= 3'b000;
				ready <= 1;
			end
		{3'b000}:
			begin
				ready <= 0;
			end
		default:
			begin
				sel <= 2'b00;
				state <= 3'b000;
				ready <= 0;
			end
		endcase
end

mux42 mux42ic0(.a(in0),.b(in168),.c(in336),.d(in504),.sel(sel),.out(mux0));
mux42 mux42ic1(.a(in1),.b(in169),.c(in337),.d(in505),.sel(sel),.out(mux1));
mux42 mux42ic2(.a(in2),.b(in170),.c(in338),.d(in506),.sel(sel),.out(mux2));
mux42 mux42ic3(.a(in3),.b(in171),.c(in339),.d(in507),.sel(sel),.out(mux3));
mux42 mux42ic4(.a(in4),.b(in172),.c(in340),.d(in508),.sel(sel),.out(mux4));
mux42 mux42ic5(.a(in5),.b(in173),.c(in341),.d(in509),.sel(sel),.out(mux5));
mux42 mux42ic6(.a(in6),.b(in174),.c(in342),.d(in510),.sel(sel),.out(mux6));
mux42 mux42ic7(.a(in7),.b(in175),.c(in343),.d(in511),.sel(sel),.out(mux7));
mux42 mux42ic8(.a(in8),.b(in176),.c(in344),.d(in512),.sel(sel),.out(mux8));
mux42 mux42ic9(.a(in9),.b(in177),.c(in345),.d(in513),.sel(sel),.out(mux9));
mux42 mux42ic10(.a(in10),.b(in178),.c(in346),.d(in514),.sel(sel),.out(mux10));
mux42 mux42ic11(.a(in11),.b(in179),.c(in347),.d(in515),.sel(sel),.out(mux11));
mux42 mux42ic12(.a(in12),.b(in180),.c(in348),.d(in516),.sel(sel),.out(mux12));
mux42 mux42ic13(.a(in13),.b(in181),.c(in349),.d(in517),.sel(sel),.out(mux13));
mux42 mux42ic14(.a(in14),.b(in182),.c(in350),.d(in518),.sel(sel),.out(mux14));
mux42 mux42ic15(.a(in15),.b(in183),.c(in351),.d(in519),.sel(sel),.out(mux15));
mux42 mux42ic16(.a(in16),.b(in184),.c(in352),.d(in520),.sel(sel),.out(mux16));
mux42 mux42ic17(.a(in17),.b(in185),.c(in353),.d(in521),.sel(sel),.out(mux17));
mux42 mux42ic18(.a(in18),.b(in186),.c(in354),.d(in522),.sel(sel),.out(mux18));
mux42 mux42ic19(.a(in19),.b(in187),.c(in355),.d(in523),.sel(sel),.out(mux19));
mux42 mux42ic20(.a(in20),.b(in188),.c(in356),.d(in524),.sel(sel),.out(mux20));
mux42 mux42ic21(.a(in21),.b(in189),.c(in357),.d(in525),.sel(sel),.out(mux21));
mux42 mux42ic22(.a(in22),.b(in190),.c(in358),.d(in526),.sel(sel),.out(mux22));
mux42 mux42ic23(.a(in23),.b(in191),.c(in359),.d(in527),.sel(sel),.out(mux23));
mux42 mux42ic24(.a(in24),.b(in192),.c(in360),.d(in528),.sel(sel),.out(mux24));
mux42 mux42ic25(.a(in25),.b(in193),.c(in361),.d(in529),.sel(sel),.out(mux25));
mux42 mux42ic26(.a(in26),.b(in194),.c(in362),.d(in530),.sel(sel),.out(mux26));
mux42 mux42ic27(.a(in27),.b(in195),.c(in363),.d(in531),.sel(sel),.out(mux27));
mux42 mux42ic28(.a(in28),.b(in196),.c(in364),.d(in532),.sel(sel),.out(mux28));
mux42 mux42ic29(.a(in29),.b(in197),.c(in365),.d(in533),.sel(sel),.out(mux29));
mux42 mux42ic30(.a(in30),.b(in198),.c(in366),.d(in534),.sel(sel),.out(mux30));
mux42 mux42ic31(.a(in31),.b(in199),.c(in367),.d(in535),.sel(sel),.out(mux31));
mux42 mux42ic32(.a(in32),.b(in200),.c(in368),.d(in536),.sel(sel),.out(mux32));
mux42 mux42ic33(.a(in33),.b(in201),.c(in369),.d(in537),.sel(sel),.out(mux33));
mux42 mux42ic34(.a(in34),.b(in202),.c(in370),.d(in538),.sel(sel),.out(mux34));
mux42 mux42ic35(.a(in35),.b(in203),.c(in371),.d(in539),.sel(sel),.out(mux35));
mux42 mux42ic36(.a(in36),.b(in204),.c(in372),.d(in540),.sel(sel),.out(mux36));
mux42 mux42ic37(.a(in37),.b(in205),.c(in373),.d(in541),.sel(sel),.out(mux37));
mux42 mux42ic38(.a(in38),.b(in206),.c(in374),.d(in542),.sel(sel),.out(mux38));
mux42 mux42ic39(.a(in39),.b(in207),.c(in375),.d(in543),.sel(sel),.out(mux39));
mux42 mux42ic40(.a(in40),.b(in208),.c(in376),.d(in544),.sel(sel),.out(mux40));
mux42 mux42ic41(.a(in41),.b(in209),.c(in377),.d(in545),.sel(sel),.out(mux41));
mux42 mux42ic42(.a(in42),.b(in210),.c(in378),.d(in546),.sel(sel),.out(mux42));
mux42 mux42ic43(.a(in43),.b(in211),.c(in379),.d(in547),.sel(sel),.out(mux43));
mux42 mux42ic44(.a(in44),.b(in212),.c(in380),.d(in548),.sel(sel),.out(mux44));
mux42 mux42ic45(.a(in45),.b(in213),.c(in381),.d(in549),.sel(sel),.out(mux45));
mux42 mux42ic46(.a(in46),.b(in214),.c(in382),.d(in550),.sel(sel),.out(mux46));
mux42 mux42ic47(.a(in47),.b(in215),.c(in383),.d(in551),.sel(sel),.out(mux47));
mux42 mux42ic48(.a(in48),.b(in216),.c(in384),.d(in552),.sel(sel),.out(mux48));
mux42 mux42ic49(.a(in49),.b(in217),.c(in385),.d(in553),.sel(sel),.out(mux49));
mux42 mux42ic50(.a(in50),.b(in218),.c(in386),.d(in554),.sel(sel),.out(mux50));
mux42 mux42ic51(.a(in51),.b(in219),.c(in387),.d(in555),.sel(sel),.out(mux51));
mux42 mux42ic52(.a(in52),.b(in220),.c(in388),.d(in556),.sel(sel),.out(mux52));
mux42 mux42ic53(.a(in53),.b(in221),.c(in389),.d(in557),.sel(sel),.out(mux53));
mux42 mux42ic54(.a(in54),.b(in222),.c(in390),.d(in558),.sel(sel),.out(mux54));
mux42 mux42ic55(.a(in55),.b(in223),.c(in391),.d(in559),.sel(sel),.out(mux55));
mux42 mux42ic56(.a(in56),.b(in224),.c(in392),.d(in560),.sel(sel),.out(mux56));
mux42 mux42ic57(.a(in57),.b(in225),.c(in393),.d(in561),.sel(sel),.out(mux57));
mux42 mux42ic58(.a(in58),.b(in226),.c(in394),.d(in562),.sel(sel),.out(mux58));
mux42 mux42ic59(.a(in59),.b(in227),.c(in395),.d(in563),.sel(sel),.out(mux59));
mux42 mux42ic60(.a(in60),.b(in228),.c(in396),.d(in564),.sel(sel),.out(mux60));
mux42 mux42ic61(.a(in61),.b(in229),.c(in397),.d(in565),.sel(sel),.out(mux61));
mux42 mux42ic62(.a(in62),.b(in230),.c(in398),.d(in566),.sel(sel),.out(mux62));
mux42 mux42ic63(.a(in63),.b(in231),.c(in399),.d(in567),.sel(sel),.out(mux63));
mux42 mux42ic64(.a(in64),.b(in232),.c(in400),.d(in568),.sel(sel),.out(mux64));
mux42 mux42ic65(.a(in65),.b(in233),.c(in401),.d(in569),.sel(sel),.out(mux65));
mux42 mux42ic66(.a(in66),.b(in234),.c(in402),.d(in570),.sel(sel),.out(mux66));
mux42 mux42ic67(.a(in67),.b(in235),.c(in403),.d(in571),.sel(sel),.out(mux67));
mux42 mux42ic68(.a(in68),.b(in236),.c(in404),.d(in572),.sel(sel),.out(mux68));
mux42 mux42ic69(.a(in69),.b(in237),.c(in405),.d(in573),.sel(sel),.out(mux69));
mux42 mux42ic70(.a(in70),.b(in238),.c(in406),.d(in574),.sel(sel),.out(mux70));
mux42 mux42ic71(.a(in71),.b(in239),.c(in407),.d(in575),.sel(sel),.out(mux71));
mux42 mux42ic72(.a(in72),.b(in240),.c(in408),.d(in576),.sel(sel),.out(mux72));
mux42 mux42ic73(.a(in73),.b(in241),.c(in409),.d(in577),.sel(sel),.out(mux73));
mux42 mux42ic74(.a(in74),.b(in242),.c(in410),.d(in578),.sel(sel),.out(mux74));
mux42 mux42ic75(.a(in75),.b(in243),.c(in411),.d(in579),.sel(sel),.out(mux75));
mux42 mux42ic76(.a(in76),.b(in244),.c(in412),.d(in580),.sel(sel),.out(mux76));
mux42 mux42ic77(.a(in77),.b(in245),.c(in413),.d(in581),.sel(sel),.out(mux77));
mux42 mux42ic78(.a(in78),.b(in246),.c(in414),.d(in582),.sel(sel),.out(mux78));
mux42 mux42ic79(.a(in79),.b(in247),.c(in415),.d(in583),.sel(sel),.out(mux79));
mux42 mux42ic80(.a(in80),.b(in248),.c(in416),.d(in584),.sel(sel),.out(mux80));
mux42 mux42ic81(.a(in81),.b(in249),.c(in417),.d(in585),.sel(sel),.out(mux81));
mux42 mux42ic82(.a(in82),.b(in250),.c(in418),.d(in586),.sel(sel),.out(mux82));
mux42 mux42ic83(.a(in83),.b(in251),.c(in419),.d(in587),.sel(sel),.out(mux83));
mux42 mux42ic84(.a(in84),.b(in252),.c(in420),.d(in588),.sel(sel),.out(mux84));
mux42 mux42ic85(.a(in85),.b(in253),.c(in421),.d(in589),.sel(sel),.out(mux85));
mux42 mux42ic86(.a(in86),.b(in254),.c(in422),.d(in590),.sel(sel),.out(mux86));
mux42 mux42ic87(.a(in87),.b(in255),.c(in423),.d(in591),.sel(sel),.out(mux87));
mux42 mux42ic88(.a(in88),.b(in256),.c(in424),.d(in592),.sel(sel),.out(mux88));
mux42 mux42ic89(.a(in89),.b(in257),.c(in425),.d(in593),.sel(sel),.out(mux89));
mux42 mux42ic90(.a(in90),.b(in258),.c(in426),.d(in594),.sel(sel),.out(mux90));
mux42 mux42ic91(.a(in91),.b(in259),.c(in427),.d(in595),.sel(sel),.out(mux91));
mux42 mux42ic92(.a(in92),.b(in260),.c(in428),.d(in596),.sel(sel),.out(mux92));
mux42 mux42ic93(.a(in93),.b(in261),.c(in429),.d(in597),.sel(sel),.out(mux93));
mux42 mux42ic94(.a(in94),.b(in262),.c(in430),.d(in598),.sel(sel),.out(mux94));
mux42 mux42ic95(.a(in95),.b(in263),.c(in431),.d(in599),.sel(sel),.out(mux95));
mux42 mux42ic96(.a(in96),.b(in264),.c(in432),.d(in600),.sel(sel),.out(mux96));
mux42 mux42ic97(.a(in97),.b(in265),.c(in433),.d(in601),.sel(sel),.out(mux97));
mux42 mux42ic98(.a(in98),.b(in266),.c(in434),.d(in602),.sel(sel),.out(mux98));
mux42 mux42ic99(.a(in99),.b(in267),.c(in435),.d(in603),.sel(sel),.out(mux99));
mux42 mux42ic100(.a(in100),.b(in268),.c(in436),.d(in604),.sel(sel),.out(mux100));
mux42 mux42ic101(.a(in101),.b(in269),.c(in437),.d(in605),.sel(sel),.out(mux101));
mux42 mux42ic102(.a(in102),.b(in270),.c(in438),.d(in606),.sel(sel),.out(mux102));
mux42 mux42ic103(.a(in103),.b(in271),.c(in439),.d(in607),.sel(sel),.out(mux103));
mux42 mux42ic104(.a(in104),.b(in272),.c(in440),.d(in608),.sel(sel),.out(mux104));
mux42 mux42ic105(.a(in105),.b(in273),.c(in441),.d(in609),.sel(sel),.out(mux105));
mux42 mux42ic106(.a(in106),.b(in274),.c(in442),.d(in610),.sel(sel),.out(mux106));
mux42 mux42ic107(.a(in107),.b(in275),.c(in443),.d(in611),.sel(sel),.out(mux107));
mux42 mux42ic108(.a(in108),.b(in276),.c(in444),.d(in612),.sel(sel),.out(mux108));
mux42 mux42ic109(.a(in109),.b(in277),.c(in445),.d(in613),.sel(sel),.out(mux109));
mux42 mux42ic110(.a(in110),.b(in278),.c(in446),.d(in614),.sel(sel),.out(mux110));
mux42 mux42ic111(.a(in111),.b(in279),.c(in447),.d(in615),.sel(sel),.out(mux111));
mux42 mux42ic112(.a(in112),.b(in280),.c(in448),.d(in616),.sel(sel),.out(mux112));
mux42 mux42ic113(.a(in113),.b(in281),.c(in449),.d(in617),.sel(sel),.out(mux113));
mux42 mux42ic114(.a(in114),.b(in282),.c(in450),.d(in618),.sel(sel),.out(mux114));
mux42 mux42ic115(.a(in115),.b(in283),.c(in451),.d(in619),.sel(sel),.out(mux115));
mux42 mux42ic116(.a(in116),.b(in284),.c(in452),.d(in620),.sel(sel),.out(mux116));
mux42 mux42ic117(.a(in117),.b(in285),.c(in453),.d(in621),.sel(sel),.out(mux117));
mux42 mux42ic118(.a(in118),.b(in286),.c(in454),.d(in622),.sel(sel),.out(mux118));
mux42 mux42ic119(.a(in119),.b(in287),.c(in455),.d(in623),.sel(sel),.out(mux119));
mux42 mux42ic120(.a(in120),.b(in288),.c(in456),.d(in624),.sel(sel),.out(mux120));
mux42 mux42ic121(.a(in121),.b(in289),.c(in457),.d(in625),.sel(sel),.out(mux121));
mux42 mux42ic122(.a(in122),.b(in290),.c(in458),.d(in626),.sel(sel),.out(mux122));
mux42 mux42ic123(.a(in123),.b(in291),.c(in459),.d(in627),.sel(sel),.out(mux123));
mux42 mux42ic124(.a(in124),.b(in292),.c(in460),.d(in628),.sel(sel),.out(mux124));
mux42 mux42ic125(.a(in125),.b(in293),.c(in461),.d(in629),.sel(sel),.out(mux125));
mux42 mux42ic126(.a(in126),.b(in294),.c(in462),.d(in630),.sel(sel),.out(mux126));
mux42 mux42ic127(.a(in127),.b(in295),.c(in463),.d(in631),.sel(sel),.out(mux127));
mux42 mux42ic128(.a(in128),.b(in296),.c(in464),.d(in632),.sel(sel),.out(mux128));
mux42 mux42ic129(.a(in129),.b(in297),.c(in465),.d(in633),.sel(sel),.out(mux129));
mux42 mux42ic130(.a(in130),.b(in298),.c(in466),.d(in634),.sel(sel),.out(mux130));
mux42 mux42ic131(.a(in131),.b(in299),.c(in467),.d(in635),.sel(sel),.out(mux131));
mux42 mux42ic132(.a(in132),.b(in300),.c(in468),.d(in636),.sel(sel),.out(mux132));
mux42 mux42ic133(.a(in133),.b(in301),.c(in469),.d(in637),.sel(sel),.out(mux133));
mux42 mux42ic134(.a(in134),.b(in302),.c(in470),.d(in638),.sel(sel),.out(mux134));
mux42 mux42ic135(.a(in135),.b(in303),.c(in471),.d(in639),.sel(sel),.out(mux135));
mux42 mux42ic136(.a(in136),.b(in304),.c(in472),.d(in640),.sel(sel),.out(mux136));
mux42 mux42ic137(.a(in137),.b(in305),.c(in473),.d(in641),.sel(sel),.out(mux137));
mux42 mux42ic138(.a(in138),.b(in306),.c(in474),.d(in642),.sel(sel),.out(mux138));
mux42 mux42ic139(.a(in139),.b(in307),.c(in475),.d(in643),.sel(sel),.out(mux139));
mux42 mux42ic140(.a(in140),.b(in308),.c(in476),.d(in644),.sel(sel),.out(mux140));
mux42 mux42ic141(.a(in141),.b(in309),.c(in477),.d(in645),.sel(sel),.out(mux141));
mux42 mux42ic142(.a(in142),.b(in310),.c(in478),.d(in646),.sel(sel),.out(mux142));
mux42 mux42ic143(.a(in143),.b(in311),.c(in479),.d(in647),.sel(sel),.out(mux143));
mux42 mux42ic144(.a(in144),.b(in312),.c(in480),.d(in648),.sel(sel),.out(mux144));
mux42 mux42ic145(.a(in145),.b(in313),.c(in481),.d(in649),.sel(sel),.out(mux145));
mux42 mux42ic146(.a(in146),.b(in314),.c(in482),.d(in650),.sel(sel),.out(mux146));
mux42 mux42ic147(.a(in147),.b(in315),.c(in483),.d(in651),.sel(sel),.out(mux147));
mux42 mux42ic148(.a(in148),.b(in316),.c(in484),.d(in652),.sel(sel),.out(mux148));
mux42 mux42ic149(.a(in149),.b(in317),.c(in485),.d(in653),.sel(sel),.out(mux149));
mux42 mux42ic150(.a(in150),.b(in318),.c(in486),.d(in654),.sel(sel),.out(mux150));
mux42 mux42ic151(.a(in151),.b(in319),.c(in487),.d(in655),.sel(sel),.out(mux151));
mux42 mux42ic152(.a(in152),.b(in320),.c(in488),.d(in656),.sel(sel),.out(mux152));
mux42 mux42ic153(.a(in153),.b(in321),.c(in489),.d(in657),.sel(sel),.out(mux153));
mux42 mux42ic154(.a(in154),.b(in322),.c(in490),.d(in658),.sel(sel),.out(mux154));
mux42 mux42ic155(.a(in155),.b(in323),.c(in491),.d(in659),.sel(sel),.out(mux155));
mux42 mux42ic156(.a(in156),.b(in324),.c(in492),.d(in660),.sel(sel),.out(mux156));
mux42 mux42ic157(.a(in157),.b(in325),.c(in493),.d(in661),.sel(sel),.out(mux157));
mux42 mux42ic158(.a(in158),.b(in326),.c(in494),.d(in662),.sel(sel),.out(mux158));
mux42 mux42ic159(.a(in159),.b(in327),.c(in495),.d(in663),.sel(sel),.out(mux159));
mux42 mux42ic160(.a(in160),.b(in328),.c(in496),.d(in664),.sel(sel),.out(mux160));
mux42 mux42ic161(.a(in161),.b(in329),.c(in497),.d(in665),.sel(sel),.out(mux161));
mux42 mux42ic162(.a(in162),.b(in330),.c(in498),.d(in666),.sel(sel),.out(mux162));
mux42 mux42ic163(.a(in163),.b(in331),.c(in499),.d(in667),.sel(sel),.out(mux163));
mux42 mux42ic164(.a(in164),.b(in332),.c(in500),.d(in668),.sel(sel),.out(mux164));
mux42 mux42ic165(.a(in165),.b(in333),.c(in501),.d(in669),.sel(sel),.out(mux165));
mux42 mux42ic166(.a(in166),.b(in334),.c(in502),.d(in670),.sel(sel),.out(mux166));
mux42 mux42ic167(.a(in167),.b(in335),.c(in503),.d(in671),.sel(sel),.out(mux167));
mux42 mux42ic168(.a(in168),.b(in336),.c(in504),.d(in672),.sel(sel),.out(mux168));
mux42 mux42ic169(.a(in169),.b(in337),.c(in505),.d(in673),.sel(sel),.out(mux169));
mux42 mux42ic170(.a(in170),.b(in338),.c(in506),.d(in674),.sel(sel),.out(mux170));
mux42 mux42ic171(.a(in171),.b(in339),.c(in507),.d(in675),.sel(sel),.out(mux171));
mux42 mux42ic172(.a(in172),.b(in340),.c(in508),.d(in676),.sel(sel),.out(mux172));
mux42 mux42ic173(.a(in173),.b(in341),.c(in509),.d(in677),.sel(sel),.out(mux173));
mux42 mux42ic174(.a(in174),.b(in342),.c(in510),.d(in678),.sel(sel),.out(mux174));
mux42 mux42ic175(.a(in175),.b(in343),.c(in511),.d(in679),.sel(sel),.out(mux175));
mux42 mux42ic176(.a(in176),.b(in344),.c(in512),.d(in680),.sel(sel),.out(mux176));
mux42 mux42ic177(.a(in177),.b(in345),.c(in513),.d(in681),.sel(sel),.out(mux177));
mux42 mux42ic178(.a(in178),.b(in346),.c(in514),.d(in682),.sel(sel),.out(mux178));
mux42 mux42ic179(.a(in179),.b(in347),.c(in515),.d(in683),.sel(sel),.out(mux179));
mux42 mux42ic180(.a(in180),.b(in348),.c(in516),.d(in684),.sel(sel),.out(mux180));
mux42 mux42ic181(.a(in181),.b(in349),.c(in517),.d(in685),.sel(sel),.out(mux181));
mux42 mux42ic182(.a(in182),.b(in350),.c(in518),.d(in686),.sel(sel),.out(mux182));
mux42 mux42ic183(.a(in183),.b(in351),.c(in519),.d(in687),.sel(sel),.out(mux183));
mux42 mux42ic184(.a(in184),.b(in352),.c(in520),.d(in688),.sel(sel),.out(mux184));
mux42 mux42ic185(.a(in185),.b(in353),.c(in521),.d(in689),.sel(sel),.out(mux185));
mux42 mux42ic186(.a(in186),.b(in354),.c(in522),.d(in690),.sel(sel),.out(mux186));
mux42 mux42ic187(.a(in187),.b(in355),.c(in523),.d(in691),.sel(sel),.out(mux187));
mux42 mux42ic188(.a(in188),.b(in356),.c(in524),.d(in692),.sel(sel),.out(mux188));
mux42 mux42ic189(.a(in189),.b(in357),.c(in525),.d(in693),.sel(sel),.out(mux189));
mux42 mux42ic190(.a(in190),.b(in358),.c(in526),.d(in694),.sel(sel),.out(mux190));
mux42 mux42ic191(.a(in191),.b(in359),.c(in527),.d(in695),.sel(sel),.out(mux191));
mux42 mux42ic192(.a(in192),.b(in360),.c(in528),.d(in696),.sel(sel),.out(mux192));
mux42 mux42ic193(.a(in193),.b(in361),.c(in529),.d(in697),.sel(sel),.out(mux193));
mux42 mux42ic194(.a(in194),.b(in362),.c(in530),.d(in698),.sel(sel),.out(mux194));
mux42 mux42ic195(.a(in195),.b(in363),.c(in531),.d(in699),.sel(sel),.out(mux195));
mux42 mux42ic196(.a(in196),.b(in364),.c(in532),.d(in700),.sel(sel),.out(mux196));
mux42 mux42ic197(.a(in197),.b(in365),.c(in533),.d(in701),.sel(sel),.out(mux197));
mux42 mux42ic198(.a(in198),.b(in366),.c(in534),.d(in702),.sel(sel),.out(mux198));
mux42 mux42ic199(.a(in199),.b(in367),.c(in535),.d(in703),.sel(sel),.out(mux199));
mux42 mux42ic200(.a(in200),.b(in368),.c(in536),.d(in704),.sel(sel),.out(mux200));
mux42 mux42ic201(.a(in201),.b(in369),.c(in537),.d(in705),.sel(sel),.out(mux201));
mux42 mux42ic202(.a(in202),.b(in370),.c(in538),.d(in706),.sel(sel),.out(mux202));
mux42 mux42ic203(.a(in203),.b(in371),.c(in539),.d(in707),.sel(sel),.out(mux203));
mux42 mux42ic204(.a(in204),.b(in372),.c(in540),.d(in708),.sel(sel),.out(mux204));
mux42 mux42ic205(.a(in205),.b(in373),.c(in541),.d(in709),.sel(sel),.out(mux205));
mux42 mux42ic206(.a(in206),.b(in374),.c(in542),.d(in710),.sel(sel),.out(mux206));
mux42 mux42ic207(.a(in207),.b(in375),.c(in543),.d(in711),.sel(sel),.out(mux207));
mux42 mux42ic208(.a(in208),.b(in376),.c(in544),.d(in712),.sel(sel),.out(mux208));
mux42 mux42ic209(.a(in209),.b(in377),.c(in545),.d(in713),.sel(sel),.out(mux209));
mux42 mux42ic210(.a(in210),.b(in378),.c(in546),.d(in714),.sel(sel),.out(mux210));
mux42 mux42ic211(.a(in211),.b(in379),.c(in547),.d(in715),.sel(sel),.out(mux211));
mux42 mux42ic212(.a(in212),.b(in380),.c(in548),.d(in716),.sel(sel),.out(mux212));
mux42 mux42ic213(.a(in213),.b(in381),.c(in549),.d(in717),.sel(sel),.out(mux213));
mux42 mux42ic214(.a(in214),.b(in382),.c(in550),.d(in718),.sel(sel),.out(mux214));
mux42 mux42ic215(.a(in215),.b(in383),.c(in551),.d(in719),.sel(sel),.out(mux215));
mux42 mux42ic216(.a(in216),.b(in384),.c(in552),.d(in720),.sel(sel),.out(mux216));
mux42 mux42ic217(.a(in217),.b(in385),.c(in553),.d(in721),.sel(sel),.out(mux217));
mux42 mux42ic218(.a(in218),.b(in386),.c(in554),.d(in722),.sel(sel),.out(mux218));
mux42 mux42ic219(.a(in219),.b(in387),.c(in555),.d(in723),.sel(sel),.out(mux219));
mux42 mux42ic220(.a(in220),.b(in388),.c(in556),.d(in724),.sel(sel),.out(mux220));
mux42 mux42ic221(.a(in221),.b(in389),.c(in557),.d(in725),.sel(sel),.out(mux221));
mux42 mux42ic222(.a(in222),.b(in390),.c(in558),.d(in726),.sel(sel),.out(mux222));
mux42 mux42ic223(.a(in223),.b(in391),.c(in559),.d(in727),.sel(sel),.out(mux223));
mux42 mux42ic224(.a(in224),.b(in392),.c(in560),.d(in728),.sel(sel),.out(mux224));
mux42 mux42ic225(.a(in225),.b(in393),.c(in561),.d(in729),.sel(sel),.out(mux225));
mux42 mux42ic226(.a(in226),.b(in394),.c(in562),.d(in730),.sel(sel),.out(mux226));
mux42 mux42ic227(.a(in227),.b(in395),.c(in563),.d(in731),.sel(sel),.out(mux227));
mux42 mux42ic228(.a(in228),.b(in396),.c(in564),.d(in732),.sel(sel),.out(mux228));
mux42 mux42ic229(.a(in229),.b(in397),.c(in565),.d(in733),.sel(sel),.out(mux229));
mux42 mux42ic230(.a(in230),.b(in398),.c(in566),.d(in734),.sel(sel),.out(mux230));
mux42 mux42ic231(.a(in231),.b(in399),.c(in567),.d(in735),.sel(sel),.out(mux231));
mux42 mux42ic232(.a(in232),.b(in400),.c(in568),.d(in736),.sel(sel),.out(mux232));
mux42 mux42ic233(.a(in233),.b(in401),.c(in569),.d(in737),.sel(sel),.out(mux233));
mux42 mux42ic234(.a(in234),.b(in402),.c(in570),.d(in738),.sel(sel),.out(mux234));
mux42 mux42ic235(.a(in235),.b(in403),.c(in571),.d(in739),.sel(sel),.out(mux235));
mux42 mux42ic236(.a(in236),.b(in404),.c(in572),.d(in740),.sel(sel),.out(mux236));
mux42 mux42ic237(.a(in237),.b(in405),.c(in573),.d(in741),.sel(sel),.out(mux237));
mux42 mux42ic238(.a(in238),.b(in406),.c(in574),.d(in742),.sel(sel),.out(mux238));
mux42 mux42ic239(.a(in239),.b(in407),.c(in575),.d(in743),.sel(sel),.out(mux239));
mux42 mux42ic240(.a(in240),.b(in408),.c(in576),.d(in744),.sel(sel),.out(mux240));
mux42 mux42ic241(.a(in241),.b(in409),.c(in577),.d(in745),.sel(sel),.out(mux241));
mux42 mux42ic242(.a(in242),.b(in410),.c(in578),.d(in746),.sel(sel),.out(mux242));
mux42 mux42ic243(.a(in243),.b(in411),.c(in579),.d(in747),.sel(sel),.out(mux243));
mux42 mux42ic244(.a(in244),.b(in412),.c(in580),.d(in748),.sel(sel),.out(mux244));
mux42 mux42ic245(.a(in245),.b(in413),.c(in581),.d(in749),.sel(sel),.out(mux245));
mux42 mux42ic246(.a(in246),.b(in414),.c(in582),.d(in750),.sel(sel),.out(mux246));
mux42 mux42ic247(.a(in247),.b(in415),.c(in583),.d(in751),.sel(sel),.out(mux247));
mux42 mux42ic248(.a(in248),.b(in416),.c(in584),.d(in752),.sel(sel),.out(mux248));
mux42 mux42ic249(.a(in249),.b(in417),.c(in585),.d(in753),.sel(sel),.out(mux249));
mux42 mux42ic250(.a(in250),.b(in418),.c(in586),.d(in754),.sel(sel),.out(mux250));
mux42 mux42ic251(.a(in251),.b(in419),.c(in587),.d(in755),.sel(sel),.out(mux251));
mux42 mux42ic252(.a(in252),.b(in420),.c(in588),.d(in756),.sel(sel),.out(mux252));
mux42 mux42ic253(.a(in253),.b(in421),.c(in589),.d(in757),.sel(sel),.out(mux253));
mux42 mux42ic254(.a(in254),.b(in422),.c(in590),.d(in758),.sel(sel),.out(mux254));
mux42 mux42ic255(.a(in255),.b(in423),.c(in591),.d(in759),.sel(sel),.out(mux255));
mux42 mux42ic256(.a(in256),.b(in424),.c(in592),.d(in760),.sel(sel),.out(mux256));
mux42 mux42ic257(.a(in257),.b(in425),.c(in593),.d(in761),.sel(sel),.out(mux257));
mux42 mux42ic258(.a(in258),.b(in426),.c(in594),.d(in762),.sel(sel),.out(mux258));
mux42 mux42ic259(.a(in259),.b(in427),.c(in595),.d(in763),.sel(sel),.out(mux259));
mux42 mux42ic260(.a(in260),.b(in428),.c(in596),.d(in764),.sel(sel),.out(mux260));
mux42 mux42ic261(.a(in261),.b(in429),.c(in597),.d(in765),.sel(sel),.out(mux261));
mux42 mux42ic262(.a(in262),.b(in430),.c(in598),.d(in766),.sel(sel),.out(mux262));
mux42 mux42ic263(.a(in263),.b(in431),.c(in599),.d(in767),.sel(sel),.out(mux263));
mux42 mux42ic264(.a(in264),.b(in432),.c(in600),.d(in768),.sel(sel),.out(mux264));
mux42 mux42ic265(.a(in265),.b(in433),.c(in601),.d(in769),.sel(sel),.out(mux265));
mux42 mux42ic266(.a(in266),.b(in434),.c(in602),.d(in770),.sel(sel),.out(mux266));
mux42 mux42ic267(.a(in267),.b(in435),.c(in603),.d(in771),.sel(sel),.out(mux267));
mux42 mux42ic268(.a(in268),.b(in436),.c(in604),.d(in772),.sel(sel),.out(mux268));
mux42 mux42ic269(.a(in269),.b(in437),.c(in605),.d(in773),.sel(sel),.out(mux269));
mux42 mux42ic270(.a(in270),.b(in438),.c(in606),.d(in774),.sel(sel),.out(mux270));
mux42 mux42ic271(.a(in271),.b(in439),.c(in607),.d(in775),.sel(sel),.out(mux271));
mux42 mux42ic272(.a(in272),.b(in440),.c(in608),.d(in776),.sel(sel),.out(mux272));
mux42 mux42ic273(.a(in273),.b(in441),.c(in609),.d(in777),.sel(sel),.out(mux273));
mux42 mux42ic274(.a(in274),.b(in442),.c(in610),.d(in778),.sel(sel),.out(mux274));
mux42 mux42ic275(.a(in275),.b(in443),.c(in611),.d(in779),.sel(sel),.out(mux275));
mux42 mux42ic276(.a(in276),.b(in444),.c(in612),.d(in780),.sel(sel),.out(mux276));
mux42 mux42ic277(.a(in277),.b(in445),.c(in613),.d(in781),.sel(sel),.out(mux277));
mux42 mux42ic278(.a(in278),.b(in446),.c(in614),.d(in782),.sel(sel),.out(mux278));
mux42 mux42ic279(.a(in279),.b(in447),.c(in615),.d(in783),.sel(sel),.out(mux279));




demux42 mux42o0(.a(conv0),.b(conv144),.c(conv288),.d(conv432),.sel(sel),.out(muxin0));
demux42 mux42o1(.a(conv1),.b(conv145),.c(conv289),.d(conv433),.sel(sel),.out(muxin1));
demux42 mux42o2(.a(conv2),.b(conv146),.c(conv290),.d(conv434),.sel(sel),.out(muxin2));
demux42 mux42o3(.a(conv3),.b(conv147),.c(conv291),.d(conv435),.sel(sel),.out(muxin3));
demux42 mux42o4(.a(conv4),.b(conv148),.c(conv292),.d(conv436),.sel(sel),.out(muxin4));
demux42 mux42o5(.a(conv5),.b(conv149),.c(conv293),.d(conv437),.sel(sel),.out(muxin5));
demux42 mux42o6(.a(conv6),.b(conv150),.c(conv294),.d(conv438),.sel(sel),.out(muxin6));
demux42 mux42o7(.a(conv7),.b(conv151),.c(conv295),.d(conv439),.sel(sel),.out(muxin7));
demux42 mux42o8(.a(conv8),.b(conv152),.c(conv296),.d(conv440),.sel(sel),.out(muxin8));
demux42 mux42o9(.a(conv9),.b(conv153),.c(conv297),.d(conv441),.sel(sel),.out(muxin9));
demux42 mux42o10(.a(conv10),.b(conv154),.c(conv298),.d(conv442),.sel(sel),.out(muxin10));
demux42 mux42o11(.a(conv11),.b(conv155),.c(conv299),.d(conv443),.sel(sel),.out(muxin11));
demux42 mux42o12(.a(conv12),.b(conv156),.c(conv300),.d(conv444),.sel(sel),.out(muxin12));
demux42 mux42o13(.a(conv13),.b(conv157),.c(conv301),.d(conv445),.sel(sel),.out(muxin13));
demux42 mux42o14(.a(conv14),.b(conv158),.c(conv302),.d(conv446),.sel(sel),.out(muxin14));
demux42 mux42o15(.a(conv15),.b(conv159),.c(conv303),.d(conv447),.sel(sel),.out(muxin15));
demux42 mux42o16(.a(conv16),.b(conv160),.c(conv304),.d(conv448),.sel(sel),.out(muxin16));
demux42 mux42o17(.a(conv17),.b(conv161),.c(conv305),.d(conv449),.sel(sel),.out(muxin17));
demux42 mux42o18(.a(conv18),.b(conv162),.c(conv306),.d(conv450),.sel(sel),.out(muxin18));
demux42 mux42o19(.a(conv19),.b(conv163),.c(conv307),.d(conv451),.sel(sel),.out(muxin19));
demux42 mux42o20(.a(conv20),.b(conv164),.c(conv308),.d(conv452),.sel(sel),.out(muxin20));
demux42 mux42o21(.a(conv21),.b(conv165),.c(conv309),.d(conv453),.sel(sel),.out(muxin21));
demux42 mux42o22(.a(conv22),.b(conv166),.c(conv310),.d(conv454),.sel(sel),.out(muxin22));
demux42 mux42o23(.a(conv23),.b(conv167),.c(conv311),.d(conv455),.sel(sel),.out(muxin23));
demux42 mux42o24(.a(conv24),.b(conv168),.c(conv312),.d(conv456),.sel(sel),.out(muxin24));
demux42 mux42o25(.a(conv25),.b(conv169),.c(conv313),.d(conv457),.sel(sel),.out(muxin25));
demux42 mux42o26(.a(conv26),.b(conv170),.c(conv314),.d(conv458),.sel(sel),.out(muxin26));
demux42 mux42o27(.a(conv27),.b(conv171),.c(conv315),.d(conv459),.sel(sel),.out(muxin27));
demux42 mux42o28(.a(conv28),.b(conv172),.c(conv316),.d(conv460),.sel(sel),.out(muxin28));
demux42 mux42o29(.a(conv29),.b(conv173),.c(conv317),.d(conv461),.sel(sel),.out(muxin29));
demux42 mux42o30(.a(conv30),.b(conv174),.c(conv318),.d(conv462),.sel(sel),.out(muxin30));
demux42 mux42o31(.a(conv31),.b(conv175),.c(conv319),.d(conv463),.sel(sel),.out(muxin31));
demux42 mux42o32(.a(conv32),.b(conv176),.c(conv320),.d(conv464),.sel(sel),.out(muxin32));
demux42 mux42o33(.a(conv33),.b(conv177),.c(conv321),.d(conv465),.sel(sel),.out(muxin33));
demux42 mux42o34(.a(conv34),.b(conv178),.c(conv322),.d(conv466),.sel(sel),.out(muxin34));
demux42 mux42o35(.a(conv35),.b(conv179),.c(conv323),.d(conv467),.sel(sel),.out(muxin35));
demux42 mux42o36(.a(conv36),.b(conv180),.c(conv324),.d(conv468),.sel(sel),.out(muxin36));
demux42 mux42o37(.a(conv37),.b(conv181),.c(conv325),.d(conv469),.sel(sel),.out(muxin37));
demux42 mux42o38(.a(conv38),.b(conv182),.c(conv326),.d(conv470),.sel(sel),.out(muxin38));
demux42 mux42o39(.a(conv39),.b(conv183),.c(conv327),.d(conv471),.sel(sel),.out(muxin39));
demux42 mux42o40(.a(conv40),.b(conv184),.c(conv328),.d(conv472),.sel(sel),.out(muxin40));
demux42 mux42o41(.a(conv41),.b(conv185),.c(conv329),.d(conv473),.sel(sel),.out(muxin41));
demux42 mux42o42(.a(conv42),.b(conv186),.c(conv330),.d(conv474),.sel(sel),.out(muxin42));
demux42 mux42o43(.a(conv43),.b(conv187),.c(conv331),.d(conv475),.sel(sel),.out(muxin43));
demux42 mux42o44(.a(conv44),.b(conv188),.c(conv332),.d(conv476),.sel(sel),.out(muxin44));
demux42 mux42o45(.a(conv45),.b(conv189),.c(conv333),.d(conv477),.sel(sel),.out(muxin45));
demux42 mux42o46(.a(conv46),.b(conv190),.c(conv334),.d(conv478),.sel(sel),.out(muxin46));
demux42 mux42o47(.a(conv47),.b(conv191),.c(conv335),.d(conv479),.sel(sel),.out(muxin47));
demux42 mux42o48(.a(conv48),.b(conv192),.c(conv336),.d(conv480),.sel(sel),.out(muxin48));
demux42 mux42o49(.a(conv49),.b(conv193),.c(conv337),.d(conv481),.sel(sel),.out(muxin49));
demux42 mux42o50(.a(conv50),.b(conv194),.c(conv338),.d(conv482),.sel(sel),.out(muxin50));
demux42 mux42o51(.a(conv51),.b(conv195),.c(conv339),.d(conv483),.sel(sel),.out(muxin51));
demux42 mux42o52(.a(conv52),.b(conv196),.c(conv340),.d(conv484),.sel(sel),.out(muxin52));
demux42 mux42o53(.a(conv53),.b(conv197),.c(conv341),.d(conv485),.sel(sel),.out(muxin53));
demux42 mux42o54(.a(conv54),.b(conv198),.c(conv342),.d(conv486),.sel(sel),.out(muxin54));
demux42 mux42o55(.a(conv55),.b(conv199),.c(conv343),.d(conv487),.sel(sel),.out(muxin55));
demux42 mux42o56(.a(conv56),.b(conv200),.c(conv344),.d(conv488),.sel(sel),.out(muxin56));
demux42 mux42o57(.a(conv57),.b(conv201),.c(conv345),.d(conv489),.sel(sel),.out(muxin57));
demux42 mux42o58(.a(conv58),.b(conv202),.c(conv346),.d(conv490),.sel(sel),.out(muxin58));
demux42 mux42o59(.a(conv59),.b(conv203),.c(conv347),.d(conv491),.sel(sel),.out(muxin59));
demux42 mux42o60(.a(conv60),.b(conv204),.c(conv348),.d(conv492),.sel(sel),.out(muxin60));
demux42 mux42o61(.a(conv61),.b(conv205),.c(conv349),.d(conv493),.sel(sel),.out(muxin61));
demux42 mux42o62(.a(conv62),.b(conv206),.c(conv350),.d(conv494),.sel(sel),.out(muxin62));
demux42 mux42o63(.a(conv63),.b(conv207),.c(conv351),.d(conv495),.sel(sel),.out(muxin63));
demux42 mux42o64(.a(conv64),.b(conv208),.c(conv352),.d(conv496),.sel(sel),.out(muxin64));
demux42 mux42o65(.a(conv65),.b(conv209),.c(conv353),.d(conv497),.sel(sel),.out(muxin65));
demux42 mux42o66(.a(conv66),.b(conv210),.c(conv354),.d(conv498),.sel(sel),.out(muxin66));
demux42 mux42o67(.a(conv67),.b(conv211),.c(conv355),.d(conv499),.sel(sel),.out(muxin67));
demux42 mux42o68(.a(conv68),.b(conv212),.c(conv356),.d(conv500),.sel(sel),.out(muxin68));
demux42 mux42o69(.a(conv69),.b(conv213),.c(conv357),.d(conv501),.sel(sel),.out(muxin69));
demux42 mux42o70(.a(conv70),.b(conv214),.c(conv358),.d(conv502),.sel(sel),.out(muxin70));
demux42 mux42o71(.a(conv71),.b(conv215),.c(conv359),.d(conv503),.sel(sel),.out(muxin71));
demux42 mux42o72(.a(conv72),.b(conv216),.c(conv360),.d(conv504),.sel(sel),.out(muxin72));
demux42 mux42o73(.a(conv73),.b(conv217),.c(conv361),.d(conv505),.sel(sel),.out(muxin73));
demux42 mux42o74(.a(conv74),.b(conv218),.c(conv362),.d(conv506),.sel(sel),.out(muxin74));
demux42 mux42o75(.a(conv75),.b(conv219),.c(conv363),.d(conv507),.sel(sel),.out(muxin75));
demux42 mux42o76(.a(conv76),.b(conv220),.c(conv364),.d(conv508),.sel(sel),.out(muxin76));
demux42 mux42o77(.a(conv77),.b(conv221),.c(conv365),.d(conv509),.sel(sel),.out(muxin77));
demux42 mux42o78(.a(conv78),.b(conv222),.c(conv366),.d(conv510),.sel(sel),.out(muxin78));
demux42 mux42o79(.a(conv79),.b(conv223),.c(conv367),.d(conv511),.sel(sel),.out(muxin79));
demux42 mux42o80(.a(conv80),.b(conv224),.c(conv368),.d(conv512),.sel(sel),.out(muxin80));
demux42 mux42o81(.a(conv81),.b(conv225),.c(conv369),.d(conv513),.sel(sel),.out(muxin81));
demux42 mux42o82(.a(conv82),.b(conv226),.c(conv370),.d(conv514),.sel(sel),.out(muxin82));
demux42 mux42o83(.a(conv83),.b(conv227),.c(conv371),.d(conv515),.sel(sel),.out(muxin83));
demux42 mux42o84(.a(conv84),.b(conv228),.c(conv372),.d(conv516),.sel(sel),.out(muxin84));
demux42 mux42o85(.a(conv85),.b(conv229),.c(conv373),.d(conv517),.sel(sel),.out(muxin85));
demux42 mux42o86(.a(conv86),.b(conv230),.c(conv374),.d(conv518),.sel(sel),.out(muxin86));
demux42 mux42o87(.a(conv87),.b(conv231),.c(conv375),.d(conv519),.sel(sel),.out(muxin87));
demux42 mux42o88(.a(conv88),.b(conv232),.c(conv376),.d(conv520),.sel(sel),.out(muxin88));
demux42 mux42o89(.a(conv89),.b(conv233),.c(conv377),.d(conv521),.sel(sel),.out(muxin89));
demux42 mux42o90(.a(conv90),.b(conv234),.c(conv378),.d(conv522),.sel(sel),.out(muxin90));
demux42 mux42o91(.a(conv91),.b(conv235),.c(conv379),.d(conv523),.sel(sel),.out(muxin91));
demux42 mux42o92(.a(conv92),.b(conv236),.c(conv380),.d(conv524),.sel(sel),.out(muxin92));
demux42 mux42o93(.a(conv93),.b(conv237),.c(conv381),.d(conv525),.sel(sel),.out(muxin93));
demux42 mux42o94(.a(conv94),.b(conv238),.c(conv382),.d(conv526),.sel(sel),.out(muxin94));
demux42 mux42o95(.a(conv95),.b(conv239),.c(conv383),.d(conv527),.sel(sel),.out(muxin95));
demux42 mux42o96(.a(conv96),.b(conv240),.c(conv384),.d(conv528),.sel(sel),.out(muxin96));
demux42 mux42o97(.a(conv97),.b(conv241),.c(conv385),.d(conv529),.sel(sel),.out(muxin97));
demux42 mux42o98(.a(conv98),.b(conv242),.c(conv386),.d(conv530),.sel(sel),.out(muxin98));
demux42 mux42o99(.a(conv99),.b(conv243),.c(conv387),.d(conv531),.sel(sel),.out(muxin99));
demux42 mux42o100(.a(conv100),.b(conv244),.c(conv388),.d(conv532),.sel(sel),.out(muxin100));
demux42 mux42o101(.a(conv101),.b(conv245),.c(conv389),.d(conv533),.sel(sel),.out(muxin101));
demux42 mux42o102(.a(conv102),.b(conv246),.c(conv390),.d(conv534),.sel(sel),.out(muxin102));
demux42 mux42o103(.a(conv103),.b(conv247),.c(conv391),.d(conv535),.sel(sel),.out(muxin103));
demux42 mux42o104(.a(conv104),.b(conv248),.c(conv392),.d(conv536),.sel(sel),.out(muxin104));
demux42 mux42o105(.a(conv105),.b(conv249),.c(conv393),.d(conv537),.sel(sel),.out(muxin105));
demux42 mux42o106(.a(conv106),.b(conv250),.c(conv394),.d(conv538),.sel(sel),.out(muxin106));
demux42 mux42o107(.a(conv107),.b(conv251),.c(conv395),.d(conv539),.sel(sel),.out(muxin107));
demux42 mux42o108(.a(conv108),.b(conv252),.c(conv396),.d(conv540),.sel(sel),.out(muxin108));
demux42 mux42o109(.a(conv109),.b(conv253),.c(conv397),.d(conv541),.sel(sel),.out(muxin109));
demux42 mux42o110(.a(conv110),.b(conv254),.c(conv398),.d(conv542),.sel(sel),.out(muxin110));
demux42 mux42o111(.a(conv111),.b(conv255),.c(conv399),.d(conv543),.sel(sel),.out(muxin111));
demux42 mux42o112(.a(conv112),.b(conv256),.c(conv400),.d(conv544),.sel(sel),.out(muxin112));
demux42 mux42o113(.a(conv113),.b(conv257),.c(conv401),.d(conv545),.sel(sel),.out(muxin113));
demux42 mux42o114(.a(conv114),.b(conv258),.c(conv402),.d(conv546),.sel(sel),.out(muxin114));
demux42 mux42o115(.a(conv115),.b(conv259),.c(conv403),.d(conv547),.sel(sel),.out(muxin115));
demux42 mux42o116(.a(conv116),.b(conv260),.c(conv404),.d(conv548),.sel(sel),.out(muxin116));
demux42 mux42o117(.a(conv117),.b(conv261),.c(conv405),.d(conv549),.sel(sel),.out(muxin117));
demux42 mux42o118(.a(conv118),.b(conv262),.c(conv406),.d(conv550),.sel(sel),.out(muxin118));
demux42 mux42o119(.a(conv119),.b(conv263),.c(conv407),.d(conv551),.sel(sel),.out(muxin119));
demux42 mux42o120(.a(conv120),.b(conv264),.c(conv408),.d(conv552),.sel(sel),.out(muxin120));
demux42 mux42o121(.a(conv121),.b(conv265),.c(conv409),.d(conv553),.sel(sel),.out(muxin121));
demux42 mux42o122(.a(conv122),.b(conv266),.c(conv410),.d(conv554),.sel(sel),.out(muxin122));
demux42 mux42o123(.a(conv123),.b(conv267),.c(conv411),.d(conv555),.sel(sel),.out(muxin123));
demux42 mux42o124(.a(conv124),.b(conv268),.c(conv412),.d(conv556),.sel(sel),.out(muxin124));
demux42 mux42o125(.a(conv125),.b(conv269),.c(conv413),.d(conv557),.sel(sel),.out(muxin125));
demux42 mux42o126(.a(conv126),.b(conv270),.c(conv414),.d(conv558),.sel(sel),.out(muxin126));
demux42 mux42o127(.a(conv127),.b(conv271),.c(conv415),.d(conv559),.sel(sel),.out(muxin127));
demux42 mux42o128(.a(conv128),.b(conv272),.c(conv416),.d(conv560),.sel(sel),.out(muxin128));
demux42 mux42o129(.a(conv129),.b(conv273),.c(conv417),.d(conv561),.sel(sel),.out(muxin129));
demux42 mux42o130(.a(conv130),.b(conv274),.c(conv418),.d(conv562),.sel(sel),.out(muxin130));
demux42 mux42o131(.a(conv131),.b(conv275),.c(conv419),.d(conv563),.sel(sel),.out(muxin131));
demux42 mux42o132(.a(conv132),.b(conv276),.c(conv420),.d(conv564),.sel(sel),.out(muxin132));
demux42 mux42o133(.a(conv133),.b(conv277),.c(conv421),.d(conv565),.sel(sel),.out(muxin133));
demux42 mux42o134(.a(conv134),.b(conv278),.c(conv422),.d(conv566),.sel(sel),.out(muxin134));
demux42 mux42o135(.a(conv135),.b(conv279),.c(conv423),.d(conv567),.sel(sel),.out(muxin135));
demux42 mux42o136(.a(conv136),.b(conv280),.c(conv424),.d(conv568),.sel(sel),.out(muxin136));
demux42 mux42o137(.a(conv137),.b(conv281),.c(conv425),.d(conv569),.sel(sel),.out(muxin137));
demux42 mux42o138(.a(conv138),.b(conv282),.c(conv426),.d(conv570),.sel(sel),.out(muxin138));
demux42 mux42o139(.a(conv139),.b(conv283),.c(conv427),.d(conv571),.sel(sel),.out(muxin139));
demux42 mux42o140(.a(conv140),.b(conv284),.c(conv428),.d(conv572),.sel(sel),.out(muxin140));
demux42 mux42o141(.a(conv141),.b(conv285),.c(conv429),.d(conv573),.sel(sel),.out(muxin141));
demux42 mux42o142(.a(conv142),.b(conv286),.c(conv430),.d(conv574),.sel(sel),.out(muxin142));
demux42 mux42o143(.a(conv143),.b(conv287),.c(conv431),.d(conv575),.sel(sel),.out(muxin143));




  Conv5D  Conv5D0(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux0),.in1(mux1),.in2(mux2),.in3(mux3),.in4(mux4),.in5(mux28),.in6(mux29),.in7(mux30),.in8(mux31),.in9(mux32),.in10(mux56),.in11(mux57),.in12(mux58),.in13(mux59),.in14(mux60),.in15(mux84),.in16(mux85),.in17(mux86),.in18(mux87),.in19(mux88),.in20(mux112),.in21(mux113),.in22(mux114),.in23(mux115),.in24(mux116), .bias(bias), .clk(clk), .out(muxin0));
 
Conv5D  Conv5D1(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux1),.in1(mux2),.in2(mux3),.in3(mux4),.in4(mux5),.in5(mux29),.in6(mux30),.in7(mux31),.in8(mux32),.in9(mux33),.in10(mux57),.in11(mux58),.in12(mux59),.in13(mux60),.in14(mux61),.in15(mux85),.in16(mux86),.in17(mux87),.in18(mux88),.in19(mux89),.in20(mux113),.in21(mux114),.in22(mux115),.in23(mux116),.in24(mux117), .bias(bias), .clk(clk), .out(muxin1));
 
Conv5D  Conv5D2(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux2),.in1(mux3),.in2(mux4),.in3(mux5),.in4(mux6),.in5(mux30),.in6(mux31),.in7(mux32),.in8(mux33),.in9(mux34),.in10(mux58),.in11(mux59),.in12(mux60),.in13(mux61),.in14(mux62),.in15(mux86),.in16(mux87),.in17(mux88),.in18(mux89),.in19(mux90),.in20(mux114),.in21(mux115),.in22(mux116),.in23(mux117),.in24(mux118), .bias(bias), .clk(clk), .out(muxin2));
 
Conv5D  Conv5D3(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux3),.in1(mux4),.in2(mux5),.in3(mux6),.in4(mux7),.in5(mux31),.in6(mux32),.in7(mux33),.in8(mux34),.in9(mux35),.in10(mux59),.in11(mux60),.in12(mux61),.in13(mux62),.in14(mux63),.in15(mux87),.in16(mux88),.in17(mux89),.in18(mux90),.in19(mux91),.in20(mux115),.in21(mux116),.in22(mux117),.in23(mux118),.in24(mux119), .bias(bias), .clk(clk), .out(muxin3));
 
Conv5D  Conv5D4(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux4),.in1(mux5),.in2(mux6),.in3(mux7),.in4(mux8),.in5(mux32),.in6(mux33),.in7(mux34),.in8(mux35),.in9(mux36),.in10(mux60),.in11(mux61),.in12(mux62),.in13(mux63),.in14(mux64),.in15(mux88),.in16(mux89),.in17(mux90),.in18(mux91),.in19(mux92),.in20(mux116),.in21(mux117),.in22(mux118),.in23(mux119),.in24(mux120), .bias(bias), .clk(clk), .out(muxin4));
 
Conv5D  Conv5D5(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux5),.in1(mux6),.in2(mux7),.in3(mux8),.in4(mux9),.in5(mux33),.in6(mux34),.in7(mux35),.in8(mux36),.in9(mux37),.in10(mux61),.in11(mux62),.in12(mux63),.in13(mux64),.in14(mux65),.in15(mux89),.in16(mux90),.in17(mux91),.in18(mux92),.in19(mux93),.in20(mux117),.in21(mux118),.in22(mux119),.in23(mux120),.in24(mux121), .bias(bias), .clk(clk), .out(muxin5));
 
Conv5D  Conv5D6(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux6),.in1(mux7),.in2(mux8),.in3(mux9),.in4(mux10),.in5(mux34),.in6(mux35),.in7(mux36),.in8(mux37),.in9(mux38),.in10(mux62),.in11(mux63),.in12(mux64),.in13(mux65),.in14(mux66),.in15(mux90),.in16(mux91),.in17(mux92),.in18(mux93),.in19(mux94),.in20(mux118),.in21(mux119),.in22(mux120),.in23(mux121),.in24(mux122), .bias(bias), .clk(clk), .out(muxin6));
 
Conv5D  Conv5D7(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux7),.in1(mux8),.in2(mux9),.in3(mux10),.in4(mux11),.in5(mux35),.in6(mux36),.in7(mux37),.in8(mux38),.in9(mux39),.in10(mux63),.in11(mux64),.in12(mux65),.in13(mux66),.in14(mux67),.in15(mux91),.in16(mux92),.in17(mux93),.in18(mux94),.in19(mux95),.in20(mux119),.in21(mux120),.in22(mux121),.in23(mux122),.in24(mux123), .bias(bias), .clk(clk), .out(muxin7));
 
Conv5D  Conv5D8(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux8),.in1(mux9),.in2(mux10),.in3(mux11),.in4(mux12),.in5(mux36),.in6(mux37),.in7(mux38),.in8(mux39),.in9(mux40),.in10(mux64),.in11(mux65),.in12(mux66),.in13(mux67),.in14(mux68),.in15(mux92),.in16(mux93),.in17(mux94),.in18(mux95),.in19(mux96),.in20(mux120),.in21(mux121),.in22(mux122),.in23(mux123),.in24(mux124), .bias(bias), .clk(clk), .out(muxin8));
 
Conv5D  Conv5D9(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux9),.in1(mux10),.in2(mux11),.in3(mux12),.in4(mux13),.in5(mux37),.in6(mux38),.in7(mux39),.in8(mux40),.in9(mux41),.in10(mux65),.in11(mux66),.in12(mux67),.in13(mux68),.in14(mux69),.in15(mux93),.in16(mux94),.in17(mux95),.in18(mux96),.in19(mux97),.in20(mux121),.in21(mux122),.in22(mux123),.in23(mux124),.in24(mux125), .bias(bias), .clk(clk), .out(muxin9));
 
Conv5D  Conv5D10(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux10),.in1(mux11),.in2(mux12),.in3(mux13),.in4(mux14),.in5(mux38),.in6(mux39),.in7(mux40),.in8(mux41),.in9(mux42),.in10(mux66),.in11(mux67),.in12(mux68),.in13(mux69),.in14(mux70),.in15(mux94),.in16(mux95),.in17(mux96),.in18(mux97),.in19(mux98),.in20(mux122),.in21(mux123),.in22(mux124),.in23(mux125),.in24(mux126), .bias(bias), .clk(clk), .out(muxin10));
 
Conv5D  Conv5D11(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux11),.in1(mux12),.in2(mux13),.in3(mux14),.in4(mux15),.in5(mux39),.in6(mux40),.in7(mux41),.in8(mux42),.in9(mux43),.in10(mux67),.in11(mux68),.in12(mux69),.in13(mux70),.in14(mux71),.in15(mux95),.in16(mux96),.in17(mux97),.in18(mux98),.in19(mux99),.in20(mux123),.in21(mux124),.in22(mux125),.in23(mux126),.in24(mux127), .bias(bias), .clk(clk), .out(muxin11));
 
Conv5D  Conv5D12(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux12),.in1(mux13),.in2(mux14),.in3(mux15),.in4(mux16),.in5(mux40),.in6(mux41),.in7(mux42),.in8(mux43),.in9(mux44),.in10(mux68),.in11(mux69),.in12(mux70),.in13(mux71),.in14(mux72),.in15(mux96),.in16(mux97),.in17(mux98),.in18(mux99),.in19(mux100),.in20(mux124),.in21(mux125),.in22(mux126),.in23(mux127),.in24(mux128), .bias(bias), .clk(clk), .out(muxin12));
 
Conv5D  Conv5D13(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux13),.in1(mux14),.in2(mux15),.in3(mux16),.in4(mux17),.in5(mux41),.in6(mux42),.in7(mux43),.in8(mux44),.in9(mux45),.in10(mux69),.in11(mux70),.in12(mux71),.in13(mux72),.in14(mux73),.in15(mux97),.in16(mux98),.in17(mux99),.in18(mux100),.in19(mux101),.in20(mux125),.in21(mux126),.in22(mux127),.in23(mux128),.in24(mux129), .bias(bias), .clk(clk), .out(muxin13));
 
Conv5D  Conv5D14(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux14),.in1(mux15),.in2(mux16),.in3(mux17),.in4(mux18),.in5(mux42),.in6(mux43),.in7(mux44),.in8(mux45),.in9(mux46),.in10(mux70),.in11(mux71),.in12(mux72),.in13(mux73),.in14(mux74),.in15(mux98),.in16(mux99),.in17(mux100),.in18(mux101),.in19(mux102),.in20(mux126),.in21(mux127),.in22(mux128),.in23(mux129),.in24(mux130), .bias(bias), .clk(clk), .out(muxin14));
 
Conv5D  Conv5D15(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux15),.in1(mux16),.in2(mux17),.in3(mux18),.in4(mux19),.in5(mux43),.in6(mux44),.in7(mux45),.in8(mux46),.in9(mux47),.in10(mux71),.in11(mux72),.in12(mux73),.in13(mux74),.in14(mux75),.in15(mux99),.in16(mux100),.in17(mux101),.in18(mux102),.in19(mux103),.in20(mux127),.in21(mux128),.in22(mux129),.in23(mux130),.in24(mux131), .bias(bias), .clk(clk), .out(muxin15));
 
Conv5D  Conv5D16(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux16),.in1(mux17),.in2(mux18),.in3(mux19),.in4(mux20),.in5(mux44),.in6(mux45),.in7(mux46),.in8(mux47),.in9(mux48),.in10(mux72),.in11(mux73),.in12(mux74),.in13(mux75),.in14(mux76),.in15(mux100),.in16(mux101),.in17(mux102),.in18(mux103),.in19(mux104),.in20(mux128),.in21(mux129),.in22(mux130),.in23(mux131),.in24(mux132), .bias(bias), .clk(clk), .out(muxin16));
 
Conv5D  Conv5D17(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux17),.in1(mux18),.in2(mux19),.in3(mux20),.in4(mux21),.in5(mux45),.in6(mux46),.in7(mux47),.in8(mux48),.in9(mux49),.in10(mux73),.in11(mux74),.in12(mux75),.in13(mux76),.in14(mux77),.in15(mux101),.in16(mux102),.in17(mux103),.in18(mux104),.in19(mux105),.in20(mux129),.in21(mux130),.in22(mux131),.in23(mux132),.in24(mux133), .bias(bias), .clk(clk), .out(muxin17));
 
Conv5D  Conv5D18(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux18),.in1(mux19),.in2(mux20),.in3(mux21),.in4(mux22),.in5(mux46),.in6(mux47),.in7(mux48),.in8(mux49),.in9(mux50),.in10(mux74),.in11(mux75),.in12(mux76),.in13(mux77),.in14(mux78),.in15(mux102),.in16(mux103),.in17(mux104),.in18(mux105),.in19(mux106),.in20(mux130),.in21(mux131),.in22(mux132),.in23(mux133),.in24(mux134), .bias(bias), .clk(clk), .out(muxin18));
 
Conv5D  Conv5D19(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux19),.in1(mux20),.in2(mux21),.in3(mux22),.in4(mux23),.in5(mux47),.in6(mux48),.in7(mux49),.in8(mux50),.in9(mux51),.in10(mux75),.in11(mux76),.in12(mux77),.in13(mux78),.in14(mux79),.in15(mux103),.in16(mux104),.in17(mux105),.in18(mux106),.in19(mux107),.in20(mux131),.in21(mux132),.in22(mux133),.in23(mux134),.in24(mux135), .bias(bias), .clk(clk), .out(muxin19));
 
Conv5D  Conv5D20(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux20),.in1(mux21),.in2(mux22),.in3(mux23),.in4(mux24),.in5(mux48),.in6(mux49),.in7(mux50),.in8(mux51),.in9(mux52),.in10(mux76),.in11(mux77),.in12(mux78),.in13(mux79),.in14(mux80),.in15(mux104),.in16(mux105),.in17(mux106),.in18(mux107),.in19(mux108),.in20(mux132),.in21(mux133),.in22(mux134),.in23(mux135),.in24(mux136), .bias(bias), .clk(clk), .out(muxin20));
 
Conv5D  Conv5D21(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux21),.in1(mux22),.in2(mux23),.in3(mux24),.in4(mux25),.in5(mux49),.in6(mux50),.in7(mux51),.in8(mux52),.in9(mux53),.in10(mux77),.in11(mux78),.in12(mux79),.in13(mux80),.in14(mux81),.in15(mux105),.in16(mux106),.in17(mux107),.in18(mux108),.in19(mux109),.in20(mux133),.in21(mux134),.in22(mux135),.in23(mux136),.in24(mux137), .bias(bias), .clk(clk), .out(muxin21));
 
Conv5D  Conv5D22(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux22),.in1(mux23),.in2(mux24),.in3(mux25),.in4(mux26),.in5(mux50),.in6(mux51),.in7(mux52),.in8(mux53),.in9(mux54),.in10(mux78),.in11(mux79),.in12(mux80),.in13(mux81),.in14(mux82),.in15(mux106),.in16(mux107),.in17(mux108),.in18(mux109),.in19(mux110),.in20(mux134),.in21(mux135),.in22(mux136),.in23(mux137),.in24(mux138), .bias(bias), .clk(clk), .out(muxin22));
 
Conv5D  Conv5D23(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux23),.in1(mux24),.in2(mux25),.in3(mux26),.in4(mux27),.in5(mux51),.in6(mux52),.in7(mux53),.in8(mux54),.in9(mux55),.in10(mux79),.in11(mux80),.in12(mux81),.in13(mux82),.in14(mux83),.in15(mux107),.in16(mux108),.in17(mux109),.in18(mux110),.in19(mux111),.in20(mux135),.in21(mux136),.in22(mux137),.in23(mux138),.in24(mux139), .bias(bias), .clk(clk), .out(muxin23));
 
Conv5D  Conv5D24(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux28),.in1(mux29),.in2(mux30),.in3(mux31),.in4(mux32),.in5(mux56),.in6(mux57),.in7(mux58),.in8(mux59),.in9(mux60),.in10(mux84),.in11(mux85),.in12(mux86),.in13(mux87),.in14(mux88),.in15(mux112),.in16(mux113),.in17(mux114),.in18(mux115),.in19(mux116),.in20(mux140),.in21(mux141),.in22(mux142),.in23(mux143),.in24(mux144), .bias(bias), .clk(clk), .out(muxin24));
 
Conv5D  Conv5D25(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux29),.in1(mux30),.in2(mux31),.in3(mux32),.in4(mux33),.in5(mux57),.in6(mux58),.in7(mux59),.in8(mux60),.in9(mux61),.in10(mux85),.in11(mux86),.in12(mux87),.in13(mux88),.in14(mux89),.in15(mux113),.in16(mux114),.in17(mux115),.in18(mux116),.in19(mux117),.in20(mux141),.in21(mux142),.in22(mux143),.in23(mux144),.in24(mux145), .bias(bias), .clk(clk), .out(muxin25));
 
Conv5D  Conv5D26(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux30),.in1(mux31),.in2(mux32),.in3(mux33),.in4(mux34),.in5(mux58),.in6(mux59),.in7(mux60),.in8(mux61),.in9(mux62),.in10(mux86),.in11(mux87),.in12(mux88),.in13(mux89),.in14(mux90),.in15(mux114),.in16(mux115),.in17(mux116),.in18(mux117),.in19(mux118),.in20(mux142),.in21(mux143),.in22(mux144),.in23(mux145),.in24(mux146), .bias(bias), .clk(clk), .out(muxin26));
 
Conv5D  Conv5D27(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux31),.in1(mux32),.in2(mux33),.in3(mux34),.in4(mux35),.in5(mux59),.in6(mux60),.in7(mux61),.in8(mux62),.in9(mux63),.in10(mux87),.in11(mux88),.in12(mux89),.in13(mux90),.in14(mux91),.in15(mux115),.in16(mux116),.in17(mux117),.in18(mux118),.in19(mux119),.in20(mux143),.in21(mux144),.in22(mux145),.in23(mux146),.in24(mux147), .bias(bias), .clk(clk), .out(muxin27));
 
Conv5D  Conv5D28(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux32),.in1(mux33),.in2(mux34),.in3(mux35),.in4(mux36),.in5(mux60),.in6(mux61),.in7(mux62),.in8(mux63),.in9(mux64),.in10(mux88),.in11(mux89),.in12(mux90),.in13(mux91),.in14(mux92),.in15(mux116),.in16(mux117),.in17(mux118),.in18(mux119),.in19(mux120),.in20(mux144),.in21(mux145),.in22(mux146),.in23(mux147),.in24(mux148), .bias(bias), .clk(clk), .out(muxin28));
 
Conv5D  Conv5D29(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux33),.in1(mux34),.in2(mux35),.in3(mux36),.in4(mux37),.in5(mux61),.in6(mux62),.in7(mux63),.in8(mux64),.in9(mux65),.in10(mux89),.in11(mux90),.in12(mux91),.in13(mux92),.in14(mux93),.in15(mux117),.in16(mux118),.in17(mux119),.in18(mux120),.in19(mux121),.in20(mux145),.in21(mux146),.in22(mux147),.in23(mux148),.in24(mux149), .bias(bias), .clk(clk), .out(muxin29));
 
Conv5D  Conv5D30(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux34),.in1(mux35),.in2(mux36),.in3(mux37),.in4(mux38),.in5(mux62),.in6(mux63),.in7(mux64),.in8(mux65),.in9(mux66),.in10(mux90),.in11(mux91),.in12(mux92),.in13(mux93),.in14(mux94),.in15(mux118),.in16(mux119),.in17(mux120),.in18(mux121),.in19(mux122),.in20(mux146),.in21(mux147),.in22(mux148),.in23(mux149),.in24(mux150), .bias(bias), .clk(clk), .out(muxin30));
 
Conv5D  Conv5D31(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux35),.in1(mux36),.in2(mux37),.in3(mux38),.in4(mux39),.in5(mux63),.in6(mux64),.in7(mux65),.in8(mux66),.in9(mux67),.in10(mux91),.in11(mux92),.in12(mux93),.in13(mux94),.in14(mux95),.in15(mux119),.in16(mux120),.in17(mux121),.in18(mux122),.in19(mux123),.in20(mux147),.in21(mux148),.in22(mux149),.in23(mux150),.in24(mux151), .bias(bias), .clk(clk), .out(muxin31));
 
Conv5D  Conv5D32(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux36),.in1(mux37),.in2(mux38),.in3(mux39),.in4(mux40),.in5(mux64),.in6(mux65),.in7(mux66),.in8(mux67),.in9(mux68),.in10(mux92),.in11(mux93),.in12(mux94),.in13(mux95),.in14(mux96),.in15(mux120),.in16(mux121),.in17(mux122),.in18(mux123),.in19(mux124),.in20(mux148),.in21(mux149),.in22(mux150),.in23(mux151),.in24(mux152), .bias(bias), .clk(clk), .out(muxin32));
 
Conv5D  Conv5D33(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux37),.in1(mux38),.in2(mux39),.in3(mux40),.in4(mux41),.in5(mux65),.in6(mux66),.in7(mux67),.in8(mux68),.in9(mux69),.in10(mux93),.in11(mux94),.in12(mux95),.in13(mux96),.in14(mux97),.in15(mux121),.in16(mux122),.in17(mux123),.in18(mux124),.in19(mux125),.in20(mux149),.in21(mux150),.in22(mux151),.in23(mux152),.in24(mux153), .bias(bias), .clk(clk), .out(muxin33));
 
Conv5D  Conv5D34(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux38),.in1(mux39),.in2(mux40),.in3(mux41),.in4(mux42),.in5(mux66),.in6(mux67),.in7(mux68),.in8(mux69),.in9(mux70),.in10(mux94),.in11(mux95),.in12(mux96),.in13(mux97),.in14(mux98),.in15(mux122),.in16(mux123),.in17(mux124),.in18(mux125),.in19(mux126),.in20(mux150),.in21(mux151),.in22(mux152),.in23(mux153),.in24(mux154), .bias(bias), .clk(clk), .out(muxin34));
 
Conv5D  Conv5D35(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux39),.in1(mux40),.in2(mux41),.in3(mux42),.in4(mux43),.in5(mux67),.in6(mux68),.in7(mux69),.in8(mux70),.in9(mux71),.in10(mux95),.in11(mux96),.in12(mux97),.in13(mux98),.in14(mux99),.in15(mux123),.in16(mux124),.in17(mux125),.in18(mux126),.in19(mux127),.in20(mux151),.in21(mux152),.in22(mux153),.in23(mux154),.in24(mux155), .bias(bias), .clk(clk), .out(muxin35));
 
Conv5D  Conv5D36(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux40),.in1(mux41),.in2(mux42),.in3(mux43),.in4(mux44),.in5(mux68),.in6(mux69),.in7(mux70),.in8(mux71),.in9(mux72),.in10(mux96),.in11(mux97),.in12(mux98),.in13(mux99),.in14(mux100),.in15(mux124),.in16(mux125),.in17(mux126),.in18(mux127),.in19(mux128),.in20(mux152),.in21(mux153),.in22(mux154),.in23(mux155),.in24(mux156), .bias(bias), .clk(clk), .out(muxin36));
 
Conv5D  Conv5D37(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux41),.in1(mux42),.in2(mux43),.in3(mux44),.in4(mux45),.in5(mux69),.in6(mux70),.in7(mux71),.in8(mux72),.in9(mux73),.in10(mux97),.in11(mux98),.in12(mux99),.in13(mux100),.in14(mux101),.in15(mux125),.in16(mux126),.in17(mux127),.in18(mux128),.in19(mux129),.in20(mux153),.in21(mux154),.in22(mux155),.in23(mux156),.in24(mux157), .bias(bias), .clk(clk), .out(muxin37));
 
Conv5D  Conv5D38(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux42),.in1(mux43),.in2(mux44),.in3(mux45),.in4(mux46),.in5(mux70),.in6(mux71),.in7(mux72),.in8(mux73),.in9(mux74),.in10(mux98),.in11(mux99),.in12(mux100),.in13(mux101),.in14(mux102),.in15(mux126),.in16(mux127),.in17(mux128),.in18(mux129),.in19(mux130),.in20(mux154),.in21(mux155),.in22(mux156),.in23(mux157),.in24(mux158), .bias(bias), .clk(clk), .out(muxin38));
 
Conv5D  Conv5D39(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux43),.in1(mux44),.in2(mux45),.in3(mux46),.in4(mux47),.in5(mux71),.in6(mux72),.in7(mux73),.in8(mux74),.in9(mux75),.in10(mux99),.in11(mux100),.in12(mux101),.in13(mux102),.in14(mux103),.in15(mux127),.in16(mux128),.in17(mux129),.in18(mux130),.in19(mux131),.in20(mux155),.in21(mux156),.in22(mux157),.in23(mux158),.in24(mux159), .bias(bias), .clk(clk), .out(muxin39));
 
Conv5D  Conv5D40(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux44),.in1(mux45),.in2(mux46),.in3(mux47),.in4(mux48),.in5(mux72),.in6(mux73),.in7(mux74),.in8(mux75),.in9(mux76),.in10(mux100),.in11(mux101),.in12(mux102),.in13(mux103),.in14(mux104),.in15(mux128),.in16(mux129),.in17(mux130),.in18(mux131),.in19(mux132),.in20(mux156),.in21(mux157),.in22(mux158),.in23(mux159),.in24(mux160), .bias(bias), .clk(clk), .out(muxin40));
 
Conv5D  Conv5D41(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux45),.in1(mux46),.in2(mux47),.in3(mux48),.in4(mux49),.in5(mux73),.in6(mux74),.in7(mux75),.in8(mux76),.in9(mux77),.in10(mux101),.in11(mux102),.in12(mux103),.in13(mux104),.in14(mux105),.in15(mux129),.in16(mux130),.in17(mux131),.in18(mux132),.in19(mux133),.in20(mux157),.in21(mux158),.in22(mux159),.in23(mux160),.in24(mux161), .bias(bias), .clk(clk), .out(muxin41));
 
Conv5D  Conv5D42(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux46),.in1(mux47),.in2(mux48),.in3(mux49),.in4(mux50),.in5(mux74),.in6(mux75),.in7(mux76),.in8(mux77),.in9(mux78),.in10(mux102),.in11(mux103),.in12(mux104),.in13(mux105),.in14(mux106),.in15(mux130),.in16(mux131),.in17(mux132),.in18(mux133),.in19(mux134),.in20(mux158),.in21(mux159),.in22(mux160),.in23(mux161),.in24(mux162), .bias(bias), .clk(clk), .out(muxin42));
 
Conv5D  Conv5D43(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux47),.in1(mux48),.in2(mux49),.in3(mux50),.in4(mux51),.in5(mux75),.in6(mux76),.in7(mux77),.in8(mux78),.in9(mux79),.in10(mux103),.in11(mux104),.in12(mux105),.in13(mux106),.in14(mux107),.in15(mux131),.in16(mux132),.in17(mux133),.in18(mux134),.in19(mux135),.in20(mux159),.in21(mux160),.in22(mux161),.in23(mux162),.in24(mux163), .bias(bias), .clk(clk), .out(muxin43));
 
Conv5D  Conv5D44(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux48),.in1(mux49),.in2(mux50),.in3(mux51),.in4(mux52),.in5(mux76),.in6(mux77),.in7(mux78),.in8(mux79),.in9(mux80),.in10(mux104),.in11(mux105),.in12(mux106),.in13(mux107),.in14(mux108),.in15(mux132),.in16(mux133),.in17(mux134),.in18(mux135),.in19(mux136),.in20(mux160),.in21(mux161),.in22(mux162),.in23(mux163),.in24(mux164), .bias(bias), .clk(clk), .out(muxin44));
 
Conv5D  Conv5D45(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux49),.in1(mux50),.in2(mux51),.in3(mux52),.in4(mux53),.in5(mux77),.in6(mux78),.in7(mux79),.in8(mux80),.in9(mux81),.in10(mux105),.in11(mux106),.in12(mux107),.in13(mux108),.in14(mux109),.in15(mux133),.in16(mux134),.in17(mux135),.in18(mux136),.in19(mux137),.in20(mux161),.in21(mux162),.in22(mux163),.in23(mux164),.in24(mux165), .bias(bias), .clk(clk), .out(muxin45));
 
Conv5D  Conv5D46(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux50),.in1(mux51),.in2(mux52),.in3(mux53),.in4(mux54),.in5(mux78),.in6(mux79),.in7(mux80),.in8(mux81),.in9(mux82),.in10(mux106),.in11(mux107),.in12(mux108),.in13(mux109),.in14(mux110),.in15(mux134),.in16(mux135),.in17(mux136),.in18(mux137),.in19(mux138),.in20(mux162),.in21(mux163),.in22(mux164),.in23(mux165),.in24(mux166), .bias(bias), .clk(clk), .out(muxin46));
 
Conv5D  Conv5D47(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux51),.in1(mux52),.in2(mux53),.in3(mux54),.in4(mux55),.in5(mux79),.in6(mux80),.in7(mux81),.in8(mux82),.in9(mux83),.in10(mux107),.in11(mux108),.in12(mux109),.in13(mux110),.in14(mux111),.in15(mux135),.in16(mux136),.in17(mux137),.in18(mux138),.in19(mux139),.in20(mux163),.in21(mux164),.in22(mux165),.in23(mux166),.in24(mux167), .bias(bias), .clk(clk), .out(muxin47));
 
Conv5D  Conv5D48(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux56),.in1(mux57),.in2(mux58),.in3(mux59),.in4(mux60),.in5(mux84),.in6(mux85),.in7(mux86),.in8(mux87),.in9(mux88),.in10(mux112),.in11(mux113),.in12(mux114),.in13(mux115),.in14(mux116),.in15(mux140),.in16(mux141),.in17(mux142),.in18(mux143),.in19(mux144),.in20(mux168),.in21(mux169),.in22(mux170),.in23(mux171),.in24(mux172), .bias(bias), .clk(clk), .out(muxin48));
 
Conv5D  Conv5D49(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux57),.in1(mux58),.in2(mux59),.in3(mux60),.in4(mux61),.in5(mux85),.in6(mux86),.in7(mux87),.in8(mux88),.in9(mux89),.in10(mux113),.in11(mux114),.in12(mux115),.in13(mux116),.in14(mux117),.in15(mux141),.in16(mux142),.in17(mux143),.in18(mux144),.in19(mux145),.in20(mux169),.in21(mux170),.in22(mux171),.in23(mux172),.in24(mux173), .bias(bias), .clk(clk), .out(muxin49));
 
Conv5D  Conv5D50(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux58),.in1(mux59),.in2(mux60),.in3(mux61),.in4(mux62),.in5(mux86),.in6(mux87),.in7(mux88),.in8(mux89),.in9(mux90),.in10(mux114),.in11(mux115),.in12(mux116),.in13(mux117),.in14(mux118),.in15(mux142),.in16(mux143),.in17(mux144),.in18(mux145),.in19(mux146),.in20(mux170),.in21(mux171),.in22(mux172),.in23(mux173),.in24(mux174), .bias(bias), .clk(clk), .out(muxin50));
 
Conv5D  Conv5D51(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux59),.in1(mux60),.in2(mux61),.in3(mux62),.in4(mux63),.in5(mux87),.in6(mux88),.in7(mux89),.in8(mux90),.in9(mux91),.in10(mux115),.in11(mux116),.in12(mux117),.in13(mux118),.in14(mux119),.in15(mux143),.in16(mux144),.in17(mux145),.in18(mux146),.in19(mux147),.in20(mux171),.in21(mux172),.in22(mux173),.in23(mux174),.in24(mux175), .bias(bias), .clk(clk), .out(muxin51));
 
Conv5D  Conv5D52(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux60),.in1(mux61),.in2(mux62),.in3(mux63),.in4(mux64),.in5(mux88),.in6(mux89),.in7(mux90),.in8(mux91),.in9(mux92),.in10(mux116),.in11(mux117),.in12(mux118),.in13(mux119),.in14(mux120),.in15(mux144),.in16(mux145),.in17(mux146),.in18(mux147),.in19(mux148),.in20(mux172),.in21(mux173),.in22(mux174),.in23(mux175),.in24(mux176), .bias(bias), .clk(clk), .out(muxin52));
 
Conv5D  Conv5D53(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux61),.in1(mux62),.in2(mux63),.in3(mux64),.in4(mux65),.in5(mux89),.in6(mux90),.in7(mux91),.in8(mux92),.in9(mux93),.in10(mux117),.in11(mux118),.in12(mux119),.in13(mux120),.in14(mux121),.in15(mux145),.in16(mux146),.in17(mux147),.in18(mux148),.in19(mux149),.in20(mux173),.in21(mux174),.in22(mux175),.in23(mux176),.in24(mux177), .bias(bias), .clk(clk), .out(muxin53));
 
Conv5D  Conv5D54(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux62),.in1(mux63),.in2(mux64),.in3(mux65),.in4(mux66),.in5(mux90),.in6(mux91),.in7(mux92),.in8(mux93),.in9(mux94),.in10(mux118),.in11(mux119),.in12(mux120),.in13(mux121),.in14(mux122),.in15(mux146),.in16(mux147),.in17(mux148),.in18(mux149),.in19(mux150),.in20(mux174),.in21(mux175),.in22(mux176),.in23(mux177),.in24(mux178), .bias(bias), .clk(clk), .out(muxin54));
 
Conv5D  Conv5D55(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux63),.in1(mux64),.in2(mux65),.in3(mux66),.in4(mux67),.in5(mux91),.in6(mux92),.in7(mux93),.in8(mux94),.in9(mux95),.in10(mux119),.in11(mux120),.in12(mux121),.in13(mux122),.in14(mux123),.in15(mux147),.in16(mux148),.in17(mux149),.in18(mux150),.in19(mux151),.in20(mux175),.in21(mux176),.in22(mux177),.in23(mux178),.in24(mux179), .bias(bias), .clk(clk), .out(muxin55));
 
Conv5D  Conv5D56(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux64),.in1(mux65),.in2(mux66),.in3(mux67),.in4(mux68),.in5(mux92),.in6(mux93),.in7(mux94),.in8(mux95),.in9(mux96),.in10(mux120),.in11(mux121),.in12(mux122),.in13(mux123),.in14(mux124),.in15(mux148),.in16(mux149),.in17(mux150),.in18(mux151),.in19(mux152),.in20(mux176),.in21(mux177),.in22(mux178),.in23(mux179),.in24(mux180), .bias(bias), .clk(clk), .out(muxin56));
 
Conv5D  Conv5D57(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux65),.in1(mux66),.in2(mux67),.in3(mux68),.in4(mux69),.in5(mux93),.in6(mux94),.in7(mux95),.in8(mux96),.in9(mux97),.in10(mux121),.in11(mux122),.in12(mux123),.in13(mux124),.in14(mux125),.in15(mux149),.in16(mux150),.in17(mux151),.in18(mux152),.in19(mux153),.in20(mux177),.in21(mux178),.in22(mux179),.in23(mux180),.in24(mux181), .bias(bias), .clk(clk), .out(muxin57));
 
Conv5D  Conv5D58(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux66),.in1(mux67),.in2(mux68),.in3(mux69),.in4(mux70),.in5(mux94),.in6(mux95),.in7(mux96),.in8(mux97),.in9(mux98),.in10(mux122),.in11(mux123),.in12(mux124),.in13(mux125),.in14(mux126),.in15(mux150),.in16(mux151),.in17(mux152),.in18(mux153),.in19(mux154),.in20(mux178),.in21(mux179),.in22(mux180),.in23(mux181),.in24(mux182), .bias(bias), .clk(clk), .out(muxin58));
 
Conv5D  Conv5D59(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux67),.in1(mux68),.in2(mux69),.in3(mux70),.in4(mux71),.in5(mux95),.in6(mux96),.in7(mux97),.in8(mux98),.in9(mux99),.in10(mux123),.in11(mux124),.in12(mux125),.in13(mux126),.in14(mux127),.in15(mux151),.in16(mux152),.in17(mux153),.in18(mux154),.in19(mux155),.in20(mux179),.in21(mux180),.in22(mux181),.in23(mux182),.in24(mux183), .bias(bias), .clk(clk), .out(muxin59));
 
Conv5D  Conv5D60(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux68),.in1(mux69),.in2(mux70),.in3(mux71),.in4(mux72),.in5(mux96),.in6(mux97),.in7(mux98),.in8(mux99),.in9(mux100),.in10(mux124),.in11(mux125),.in12(mux126),.in13(mux127),.in14(mux128),.in15(mux152),.in16(mux153),.in17(mux154),.in18(mux155),.in19(mux156),.in20(mux180),.in21(mux181),.in22(mux182),.in23(mux183),.in24(mux184), .bias(bias), .clk(clk), .out(muxin60));
 
Conv5D  Conv5D61(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux69),.in1(mux70),.in2(mux71),.in3(mux72),.in4(mux73),.in5(mux97),.in6(mux98),.in7(mux99),.in8(mux100),.in9(mux101),.in10(mux125),.in11(mux126),.in12(mux127),.in13(mux128),.in14(mux129),.in15(mux153),.in16(mux154),.in17(mux155),.in18(mux156),.in19(mux157),.in20(mux181),.in21(mux182),.in22(mux183),.in23(mux184),.in24(mux185), .bias(bias), .clk(clk), .out(muxin61));
 
Conv5D  Conv5D62(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux70),.in1(mux71),.in2(mux72),.in3(mux73),.in4(mux74),.in5(mux98),.in6(mux99),.in7(mux100),.in8(mux101),.in9(mux102),.in10(mux126),.in11(mux127),.in12(mux128),.in13(mux129),.in14(mux130),.in15(mux154),.in16(mux155),.in17(mux156),.in18(mux157),.in19(mux158),.in20(mux182),.in21(mux183),.in22(mux184),.in23(mux185),.in24(mux186), .bias(bias), .clk(clk), .out(muxin62));
 
Conv5D  Conv5D63(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux71),.in1(mux72),.in2(mux73),.in3(mux74),.in4(mux75),.in5(mux99),.in6(mux100),.in7(mux101),.in8(mux102),.in9(mux103),.in10(mux127),.in11(mux128),.in12(mux129),.in13(mux130),.in14(mux131),.in15(mux155),.in16(mux156),.in17(mux157),.in18(mux158),.in19(mux159),.in20(mux183),.in21(mux184),.in22(mux185),.in23(mux186),.in24(mux187), .bias(bias), .clk(clk), .out(muxin63));
 
Conv5D  Conv5D64(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux72),.in1(mux73),.in2(mux74),.in3(mux75),.in4(mux76),.in5(mux100),.in6(mux101),.in7(mux102),.in8(mux103),.in9(mux104),.in10(mux128),.in11(mux129),.in12(mux130),.in13(mux131),.in14(mux132),.in15(mux156),.in16(mux157),.in17(mux158),.in18(mux159),.in19(mux160),.in20(mux184),.in21(mux185),.in22(mux186),.in23(mux187),.in24(mux188), .bias(bias), .clk(clk), .out(muxin64));
 
Conv5D  Conv5D65(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux73),.in1(mux74),.in2(mux75),.in3(mux76),.in4(mux77),.in5(mux101),.in6(mux102),.in7(mux103),.in8(mux104),.in9(mux105),.in10(mux129),.in11(mux130),.in12(mux131),.in13(mux132),.in14(mux133),.in15(mux157),.in16(mux158),.in17(mux159),.in18(mux160),.in19(mux161),.in20(mux185),.in21(mux186),.in22(mux187),.in23(mux188),.in24(mux189), .bias(bias), .clk(clk), .out(muxin65));
 
Conv5D  Conv5D66(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux74),.in1(mux75),.in2(mux76),.in3(mux77),.in4(mux78),.in5(mux102),.in6(mux103),.in7(mux104),.in8(mux105),.in9(mux106),.in10(mux130),.in11(mux131),.in12(mux132),.in13(mux133),.in14(mux134),.in15(mux158),.in16(mux159),.in17(mux160),.in18(mux161),.in19(mux162),.in20(mux186),.in21(mux187),.in22(mux188),.in23(mux189),.in24(mux190), .bias(bias), .clk(clk), .out(muxin66));
 
Conv5D  Conv5D67(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux75),.in1(mux76),.in2(mux77),.in3(mux78),.in4(mux79),.in5(mux103),.in6(mux104),.in7(mux105),.in8(mux106),.in9(mux107),.in10(mux131),.in11(mux132),.in12(mux133),.in13(mux134),.in14(mux135),.in15(mux159),.in16(mux160),.in17(mux161),.in18(mux162),.in19(mux163),.in20(mux187),.in21(mux188),.in22(mux189),.in23(mux190),.in24(mux191), .bias(bias), .clk(clk), .out(muxin67));
 
Conv5D  Conv5D68(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux76),.in1(mux77),.in2(mux78),.in3(mux79),.in4(mux80),.in5(mux104),.in6(mux105),.in7(mux106),.in8(mux107),.in9(mux108),.in10(mux132),.in11(mux133),.in12(mux134),.in13(mux135),.in14(mux136),.in15(mux160),.in16(mux161),.in17(mux162),.in18(mux163),.in19(mux164),.in20(mux188),.in21(mux189),.in22(mux190),.in23(mux191),.in24(mux192), .bias(bias), .clk(clk), .out(muxin68));
 
Conv5D  Conv5D69(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux77),.in1(mux78),.in2(mux79),.in3(mux80),.in4(mux81),.in5(mux105),.in6(mux106),.in7(mux107),.in8(mux108),.in9(mux109),.in10(mux133),.in11(mux134),.in12(mux135),.in13(mux136),.in14(mux137),.in15(mux161),.in16(mux162),.in17(mux163),.in18(mux164),.in19(mux165),.in20(mux189),.in21(mux190),.in22(mux191),.in23(mux192),.in24(mux193), .bias(bias), .clk(clk), .out(muxin69));
 
Conv5D  Conv5D70(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux78),.in1(mux79),.in2(mux80),.in3(mux81),.in4(mux82),.in5(mux106),.in6(mux107),.in7(mux108),.in8(mux109),.in9(mux110),.in10(mux134),.in11(mux135),.in12(mux136),.in13(mux137),.in14(mux138),.in15(mux162),.in16(mux163),.in17(mux164),.in18(mux165),.in19(mux166),.in20(mux190),.in21(mux191),.in22(mux192),.in23(mux193),.in24(mux194), .bias(bias), .clk(clk), .out(muxin70));
 
Conv5D  Conv5D71(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux79),.in1(mux80),.in2(mux81),.in3(mux82),.in4(mux83),.in5(mux107),.in6(mux108),.in7(mux109),.in8(mux110),.in9(mux111),.in10(mux135),.in11(mux136),.in12(mux137),.in13(mux138),.in14(mux139),.in15(mux163),.in16(mux164),.in17(mux165),.in18(mux166),.in19(mux167),.in20(mux191),.in21(mux192),.in22(mux193),.in23(mux194),.in24(mux195), .bias(bias), .clk(clk), .out(muxin71));
 
Conv5D  Conv5D72(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux84),.in1(mux85),.in2(mux86),.in3(mux87),.in4(mux88),.in5(mux112),.in6(mux113),.in7(mux114),.in8(mux115),.in9(mux116),.in10(mux140),.in11(mux141),.in12(mux142),.in13(mux143),.in14(mux144),.in15(mux168),.in16(mux169),.in17(mux170),.in18(mux171),.in19(mux172),.in20(mux196),.in21(mux197),.in22(mux198),.in23(mux199),.in24(mux200), .bias(bias), .clk(clk), .out(muxin72));
 
Conv5D  Conv5D73(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux85),.in1(mux86),.in2(mux87),.in3(mux88),.in4(mux89),.in5(mux113),.in6(mux114),.in7(mux115),.in8(mux116),.in9(mux117),.in10(mux141),.in11(mux142),.in12(mux143),.in13(mux144),.in14(mux145),.in15(mux169),.in16(mux170),.in17(mux171),.in18(mux172),.in19(mux173),.in20(mux197),.in21(mux198),.in22(mux199),.in23(mux200),.in24(mux201), .bias(bias), .clk(clk), .out(muxin73));
 
Conv5D  Conv5D74(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux86),.in1(mux87),.in2(mux88),.in3(mux89),.in4(mux90),.in5(mux114),.in6(mux115),.in7(mux116),.in8(mux117),.in9(mux118),.in10(mux142),.in11(mux143),.in12(mux144),.in13(mux145),.in14(mux146),.in15(mux170),.in16(mux171),.in17(mux172),.in18(mux173),.in19(mux174),.in20(mux198),.in21(mux199),.in22(mux200),.in23(mux201),.in24(mux202), .bias(bias), .clk(clk), .out(muxin74));
 
Conv5D  Conv5D75(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux87),.in1(mux88),.in2(mux89),.in3(mux90),.in4(mux91),.in5(mux115),.in6(mux116),.in7(mux117),.in8(mux118),.in9(mux119),.in10(mux143),.in11(mux144),.in12(mux145),.in13(mux146),.in14(mux147),.in15(mux171),.in16(mux172),.in17(mux173),.in18(mux174),.in19(mux175),.in20(mux199),.in21(mux200),.in22(mux201),.in23(mux202),.in24(mux203), .bias(bias), .clk(clk), .out(muxin75));
 
Conv5D  Conv5D76(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux88),.in1(mux89),.in2(mux90),.in3(mux91),.in4(mux92),.in5(mux116),.in6(mux117),.in7(mux118),.in8(mux119),.in9(mux120),.in10(mux144),.in11(mux145),.in12(mux146),.in13(mux147),.in14(mux148),.in15(mux172),.in16(mux173),.in17(mux174),.in18(mux175),.in19(mux176),.in20(mux200),.in21(mux201),.in22(mux202),.in23(mux203),.in24(mux204), .bias(bias), .clk(clk), .out(muxin76));
 
Conv5D  Conv5D77(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux89),.in1(mux90),.in2(mux91),.in3(mux92),.in4(mux93),.in5(mux117),.in6(mux118),.in7(mux119),.in8(mux120),.in9(mux121),.in10(mux145),.in11(mux146),.in12(mux147),.in13(mux148),.in14(mux149),.in15(mux173),.in16(mux174),.in17(mux175),.in18(mux176),.in19(mux177),.in20(mux201),.in21(mux202),.in22(mux203),.in23(mux204),.in24(mux205), .bias(bias), .clk(clk), .out(muxin77));
 
Conv5D  Conv5D78(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux90),.in1(mux91),.in2(mux92),.in3(mux93),.in4(mux94),.in5(mux118),.in6(mux119),.in7(mux120),.in8(mux121),.in9(mux122),.in10(mux146),.in11(mux147),.in12(mux148),.in13(mux149),.in14(mux150),.in15(mux174),.in16(mux175),.in17(mux176),.in18(mux177),.in19(mux178),.in20(mux202),.in21(mux203),.in22(mux204),.in23(mux205),.in24(mux206), .bias(bias), .clk(clk), .out(muxin78));
 
Conv5D  Conv5D79(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux91),.in1(mux92),.in2(mux93),.in3(mux94),.in4(mux95),.in5(mux119),.in6(mux120),.in7(mux121),.in8(mux122),.in9(mux123),.in10(mux147),.in11(mux148),.in12(mux149),.in13(mux150),.in14(mux151),.in15(mux175),.in16(mux176),.in17(mux177),.in18(mux178),.in19(mux179),.in20(mux203),.in21(mux204),.in22(mux205),.in23(mux206),.in24(mux207), .bias(bias), .clk(clk), .out(muxin79));
 
Conv5D  Conv5D80(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux92),.in1(mux93),.in2(mux94),.in3(mux95),.in4(mux96),.in5(mux120),.in6(mux121),.in7(mux122),.in8(mux123),.in9(mux124),.in10(mux148),.in11(mux149),.in12(mux150),.in13(mux151),.in14(mux152),.in15(mux176),.in16(mux177),.in17(mux178),.in18(mux179),.in19(mux180),.in20(mux204),.in21(mux205),.in22(mux206),.in23(mux207),.in24(mux208), .bias(bias), .clk(clk), .out(muxin80));
 
Conv5D  Conv5D81(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux93),.in1(mux94),.in2(mux95),.in3(mux96),.in4(mux97),.in5(mux121),.in6(mux122),.in7(mux123),.in8(mux124),.in9(mux125),.in10(mux149),.in11(mux150),.in12(mux151),.in13(mux152),.in14(mux153),.in15(mux177),.in16(mux178),.in17(mux179),.in18(mux180),.in19(mux181),.in20(mux205),.in21(mux206),.in22(mux207),.in23(mux208),.in24(mux209), .bias(bias), .clk(clk), .out(muxin81));
 
Conv5D  Conv5D82(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux94),.in1(mux95),.in2(mux96),.in3(mux97),.in4(mux98),.in5(mux122),.in6(mux123),.in7(mux124),.in8(mux125),.in9(mux126),.in10(mux150),.in11(mux151),.in12(mux152),.in13(mux153),.in14(mux154),.in15(mux178),.in16(mux179),.in17(mux180),.in18(mux181),.in19(mux182),.in20(mux206),.in21(mux207),.in22(mux208),.in23(mux209),.in24(mux210), .bias(bias), .clk(clk), .out(muxin82));
 
Conv5D  Conv5D83(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux95),.in1(mux96),.in2(mux97),.in3(mux98),.in4(mux99),.in5(mux123),.in6(mux124),.in7(mux125),.in8(mux126),.in9(mux127),.in10(mux151),.in11(mux152),.in12(mux153),.in13(mux154),.in14(mux155),.in15(mux179),.in16(mux180),.in17(mux181),.in18(mux182),.in19(mux183),.in20(mux207),.in21(mux208),.in22(mux209),.in23(mux210),.in24(mux211), .bias(bias), .clk(clk), .out(muxin83));
 
Conv5D  Conv5D84(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux96),.in1(mux97),.in2(mux98),.in3(mux99),.in4(mux100),.in5(mux124),.in6(mux125),.in7(mux126),.in8(mux127),.in9(mux128),.in10(mux152),.in11(mux153),.in12(mux154),.in13(mux155),.in14(mux156),.in15(mux180),.in16(mux181),.in17(mux182),.in18(mux183),.in19(mux184),.in20(mux208),.in21(mux209),.in22(mux210),.in23(mux211),.in24(mux212), .bias(bias), .clk(clk), .out(muxin84));
 
Conv5D  Conv5D85(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux97),.in1(mux98),.in2(mux99),.in3(mux100),.in4(mux101),.in5(mux125),.in6(mux126),.in7(mux127),.in8(mux128),.in9(mux129),.in10(mux153),.in11(mux154),.in12(mux155),.in13(mux156),.in14(mux157),.in15(mux181),.in16(mux182),.in17(mux183),.in18(mux184),.in19(mux185),.in20(mux209),.in21(mux210),.in22(mux211),.in23(mux212),.in24(mux213), .bias(bias), .clk(clk), .out(muxin85));
 
Conv5D  Conv5D86(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux98),.in1(mux99),.in2(mux100),.in3(mux101),.in4(mux102),.in5(mux126),.in6(mux127),.in7(mux128),.in8(mux129),.in9(mux130),.in10(mux154),.in11(mux155),.in12(mux156),.in13(mux157),.in14(mux158),.in15(mux182),.in16(mux183),.in17(mux184),.in18(mux185),.in19(mux186),.in20(mux210),.in21(mux211),.in22(mux212),.in23(mux213),.in24(mux214), .bias(bias), .clk(clk), .out(muxin86));
 
Conv5D  Conv5D87(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux99),.in1(mux100),.in2(mux101),.in3(mux102),.in4(mux103),.in5(mux127),.in6(mux128),.in7(mux129),.in8(mux130),.in9(mux131),.in10(mux155),.in11(mux156),.in12(mux157),.in13(mux158),.in14(mux159),.in15(mux183),.in16(mux184),.in17(mux185),.in18(mux186),.in19(mux187),.in20(mux211),.in21(mux212),.in22(mux213),.in23(mux214),.in24(mux215), .bias(bias), .clk(clk), .out(muxin87));
 
Conv5D  Conv5D88(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux100),.in1(mux101),.in2(mux102),.in3(mux103),.in4(mux104),.in5(mux128),.in6(mux129),.in7(mux130),.in8(mux131),.in9(mux132),.in10(mux156),.in11(mux157),.in12(mux158),.in13(mux159),.in14(mux160),.in15(mux184),.in16(mux185),.in17(mux186),.in18(mux187),.in19(mux188),.in20(mux212),.in21(mux213),.in22(mux214),.in23(mux215),.in24(mux216), .bias(bias), .clk(clk), .out(muxin88));
 
Conv5D  Conv5D89(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux101),.in1(mux102),.in2(mux103),.in3(mux104),.in4(mux105),.in5(mux129),.in6(mux130),.in7(mux131),.in8(mux132),.in9(mux133),.in10(mux157),.in11(mux158),.in12(mux159),.in13(mux160),.in14(mux161),.in15(mux185),.in16(mux186),.in17(mux187),.in18(mux188),.in19(mux189),.in20(mux213),.in21(mux214),.in22(mux215),.in23(mux216),.in24(mux217), .bias(bias), .clk(clk), .out(muxin89));
 
Conv5D  Conv5D90(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux102),.in1(mux103),.in2(mux104),.in3(mux105),.in4(mux106),.in5(mux130),.in6(mux131),.in7(mux132),.in8(mux133),.in9(mux134),.in10(mux158),.in11(mux159),.in12(mux160),.in13(mux161),.in14(mux162),.in15(mux186),.in16(mux187),.in17(mux188),.in18(mux189),.in19(mux190),.in20(mux214),.in21(mux215),.in22(mux216),.in23(mux217),.in24(mux218), .bias(bias), .clk(clk), .out(muxin90));
 
Conv5D  Conv5D91(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux103),.in1(mux104),.in2(mux105),.in3(mux106),.in4(mux107),.in5(mux131),.in6(mux132),.in7(mux133),.in8(mux134),.in9(mux135),.in10(mux159),.in11(mux160),.in12(mux161),.in13(mux162),.in14(mux163),.in15(mux187),.in16(mux188),.in17(mux189),.in18(mux190),.in19(mux191),.in20(mux215),.in21(mux216),.in22(mux217),.in23(mux218),.in24(mux219), .bias(bias), .clk(clk), .out(muxin91));
 
Conv5D  Conv5D92(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux104),.in1(mux105),.in2(mux106),.in3(mux107),.in4(mux108),.in5(mux132),.in6(mux133),.in7(mux134),.in8(mux135),.in9(mux136),.in10(mux160),.in11(mux161),.in12(mux162),.in13(mux163),.in14(mux164),.in15(mux188),.in16(mux189),.in17(mux190),.in18(mux191),.in19(mux192),.in20(mux216),.in21(mux217),.in22(mux218),.in23(mux219),.in24(mux220), .bias(bias), .clk(clk), .out(muxin92));
 
Conv5D  Conv5D93(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux105),.in1(mux106),.in2(mux107),.in3(mux108),.in4(mux109),.in5(mux133),.in6(mux134),.in7(mux135),.in8(mux136),.in9(mux137),.in10(mux161),.in11(mux162),.in12(mux163),.in13(mux164),.in14(mux165),.in15(mux189),.in16(mux190),.in17(mux191),.in18(mux192),.in19(mux193),.in20(mux217),.in21(mux218),.in22(mux219),.in23(mux220),.in24(mux221), .bias(bias), .clk(clk), .out(muxin93));
 
Conv5D  Conv5D94(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux106),.in1(mux107),.in2(mux108),.in3(mux109),.in4(mux110),.in5(mux134),.in6(mux135),.in7(mux136),.in8(mux137),.in9(mux138),.in10(mux162),.in11(mux163),.in12(mux164),.in13(mux165),.in14(mux166),.in15(mux190),.in16(mux191),.in17(mux192),.in18(mux193),.in19(mux194),.in20(mux218),.in21(mux219),.in22(mux220),.in23(mux221),.in24(mux222), .bias(bias), .clk(clk), .out(muxin94));
 
Conv5D  Conv5D95(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux107),.in1(mux108),.in2(mux109),.in3(mux110),.in4(mux111),.in5(mux135),.in6(mux136),.in7(mux137),.in8(mux138),.in9(mux139),.in10(mux163),.in11(mux164),.in12(mux165),.in13(mux166),.in14(mux167),.in15(mux191),.in16(mux192),.in17(mux193),.in18(mux194),.in19(mux195),.in20(mux219),.in21(mux220),.in22(mux221),.in23(mux222),.in24(mux223), .bias(bias), .clk(clk), .out(muxin95));
 
Conv5D  Conv5D96(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux112),.in1(mux113),.in2(mux114),.in3(mux115),.in4(mux116),.in5(mux140),.in6(mux141),.in7(mux142),.in8(mux143),.in9(mux144),.in10(mux168),.in11(mux169),.in12(mux170),.in13(mux171),.in14(mux172),.in15(mux196),.in16(mux197),.in17(mux198),.in18(mux199),.in19(mux200),.in20(mux224),.in21(mux225),.in22(mux226),.in23(mux227),.in24(mux228), .bias(bias), .clk(clk), .out(muxin96));
 
Conv5D  Conv5D97(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux113),.in1(mux114),.in2(mux115),.in3(mux116),.in4(mux117),.in5(mux141),.in6(mux142),.in7(mux143),.in8(mux144),.in9(mux145),.in10(mux169),.in11(mux170),.in12(mux171),.in13(mux172),.in14(mux173),.in15(mux197),.in16(mux198),.in17(mux199),.in18(mux200),.in19(mux201),.in20(mux225),.in21(mux226),.in22(mux227),.in23(mux228),.in24(mux229), .bias(bias), .clk(clk), .out(muxin97));
 
Conv5D  Conv5D98(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux114),.in1(mux115),.in2(mux116),.in3(mux117),.in4(mux118),.in5(mux142),.in6(mux143),.in7(mux144),.in8(mux145),.in9(mux146),.in10(mux170),.in11(mux171),.in12(mux172),.in13(mux173),.in14(mux174),.in15(mux198),.in16(mux199),.in17(mux200),.in18(mux201),.in19(mux202),.in20(mux226),.in21(mux227),.in22(mux228),.in23(mux229),.in24(mux230), .bias(bias), .clk(clk), .out(muxin98));
 
Conv5D  Conv5D99(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux115),.in1(mux116),.in2(mux117),.in3(mux118),.in4(mux119),.in5(mux143),.in6(mux144),.in7(mux145),.in8(mux146),.in9(mux147),.in10(mux171),.in11(mux172),.in12(mux173),.in13(mux174),.in14(mux175),.in15(mux199),.in16(mux200),.in17(mux201),.in18(mux202),.in19(mux203),.in20(mux227),.in21(mux228),.in22(mux229),.in23(mux230),.in24(mux231), .bias(bias), .clk(clk), .out(muxin99));
 
Conv5D  Conv5D100(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux116),.in1(mux117),.in2(mux118),.in3(mux119),.in4(mux120),.in5(mux144),.in6(mux145),.in7(mux146),.in8(mux147),.in9(mux148),.in10(mux172),.in11(mux173),.in12(mux174),.in13(mux175),.in14(mux176),.in15(mux200),.in16(mux201),.in17(mux202),.in18(mux203),.in19(mux204),.in20(mux228),.in21(mux229),.in22(mux230),.in23(mux231),.in24(mux232), .bias(bias), .clk(clk), .out(muxin100));
 
Conv5D  Conv5D101(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux117),.in1(mux118),.in2(mux119),.in3(mux120),.in4(mux121),.in5(mux145),.in6(mux146),.in7(mux147),.in8(mux148),.in9(mux149),.in10(mux173),.in11(mux174),.in12(mux175),.in13(mux176),.in14(mux177),.in15(mux201),.in16(mux202),.in17(mux203),.in18(mux204),.in19(mux205),.in20(mux229),.in21(mux230),.in22(mux231),.in23(mux232),.in24(mux233), .bias(bias), .clk(clk), .out(muxin101));
 
Conv5D  Conv5D102(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux118),.in1(mux119),.in2(mux120),.in3(mux121),.in4(mux122),.in5(mux146),.in6(mux147),.in7(mux148),.in8(mux149),.in9(mux150),.in10(mux174),.in11(mux175),.in12(mux176),.in13(mux177),.in14(mux178),.in15(mux202),.in16(mux203),.in17(mux204),.in18(mux205),.in19(mux206),.in20(mux230),.in21(mux231),.in22(mux232),.in23(mux233),.in24(mux234), .bias(bias), .clk(clk), .out(muxin102));
 
Conv5D  Conv5D103(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux119),.in1(mux120),.in2(mux121),.in3(mux122),.in4(mux123),.in5(mux147),.in6(mux148),.in7(mux149),.in8(mux150),.in9(mux151),.in10(mux175),.in11(mux176),.in12(mux177),.in13(mux178),.in14(mux179),.in15(mux203),.in16(mux204),.in17(mux205),.in18(mux206),.in19(mux207),.in20(mux231),.in21(mux232),.in22(mux233),.in23(mux234),.in24(mux235), .bias(bias), .clk(clk), .out(muxin103));
 
Conv5D  Conv5D104(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux120),.in1(mux121),.in2(mux122),.in3(mux123),.in4(mux124),.in5(mux148),.in6(mux149),.in7(mux150),.in8(mux151),.in9(mux152),.in10(mux176),.in11(mux177),.in12(mux178),.in13(mux179),.in14(mux180),.in15(mux204),.in16(mux205),.in17(mux206),.in18(mux207),.in19(mux208),.in20(mux232),.in21(mux233),.in22(mux234),.in23(mux235),.in24(mux236), .bias(bias), .clk(clk), .out(muxin104));
 
Conv5D  Conv5D105(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux121),.in1(mux122),.in2(mux123),.in3(mux124),.in4(mux125),.in5(mux149),.in6(mux150),.in7(mux151),.in8(mux152),.in9(mux153),.in10(mux177),.in11(mux178),.in12(mux179),.in13(mux180),.in14(mux181),.in15(mux205),.in16(mux206),.in17(mux207),.in18(mux208),.in19(mux209),.in20(mux233),.in21(mux234),.in22(mux235),.in23(mux236),.in24(mux237), .bias(bias), .clk(clk), .out(muxin105));
 
Conv5D  Conv5D106(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux122),.in1(mux123),.in2(mux124),.in3(mux125),.in4(mux126),.in5(mux150),.in6(mux151),.in7(mux152),.in8(mux153),.in9(mux154),.in10(mux178),.in11(mux179),.in12(mux180),.in13(mux181),.in14(mux182),.in15(mux206),.in16(mux207),.in17(mux208),.in18(mux209),.in19(mux210),.in20(mux234),.in21(mux235),.in22(mux236),.in23(mux237),.in24(mux238), .bias(bias), .clk(clk), .out(muxin106));
 
Conv5D  Conv5D107(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux123),.in1(mux124),.in2(mux125),.in3(mux126),.in4(mux127),.in5(mux151),.in6(mux152),.in7(mux153),.in8(mux154),.in9(mux155),.in10(mux179),.in11(mux180),.in12(mux181),.in13(mux182),.in14(mux183),.in15(mux207),.in16(mux208),.in17(mux209),.in18(mux210),.in19(mux211),.in20(mux235),.in21(mux236),.in22(mux237),.in23(mux238),.in24(mux239), .bias(bias), .clk(clk), .out(muxin107));
 
Conv5D  Conv5D108(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux124),.in1(mux125),.in2(mux126),.in3(mux127),.in4(mux128),.in5(mux152),.in6(mux153),.in7(mux154),.in8(mux155),.in9(mux156),.in10(mux180),.in11(mux181),.in12(mux182),.in13(mux183),.in14(mux184),.in15(mux208),.in16(mux209),.in17(mux210),.in18(mux211),.in19(mux212),.in20(mux236),.in21(mux237),.in22(mux238),.in23(mux239),.in24(mux240), .bias(bias), .clk(clk), .out(muxin108));
 
Conv5D  Conv5D109(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux125),.in1(mux126),.in2(mux127),.in3(mux128),.in4(mux129),.in5(mux153),.in6(mux154),.in7(mux155),.in8(mux156),.in9(mux157),.in10(mux181),.in11(mux182),.in12(mux183),.in13(mux184),.in14(mux185),.in15(mux209),.in16(mux210),.in17(mux211),.in18(mux212),.in19(mux213),.in20(mux237),.in21(mux238),.in22(mux239),.in23(mux240),.in24(mux241), .bias(bias), .clk(clk), .out(muxin109));
 
Conv5D  Conv5D110(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux126),.in1(mux127),.in2(mux128),.in3(mux129),.in4(mux130),.in5(mux154),.in6(mux155),.in7(mux156),.in8(mux157),.in9(mux158),.in10(mux182),.in11(mux183),.in12(mux184),.in13(mux185),.in14(mux186),.in15(mux210),.in16(mux211),.in17(mux212),.in18(mux213),.in19(mux214),.in20(mux238),.in21(mux239),.in22(mux240),.in23(mux241),.in24(mux242), .bias(bias), .clk(clk), .out(muxin110));
 
Conv5D  Conv5D111(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux127),.in1(mux128),.in2(mux129),.in3(mux130),.in4(mux131),.in5(mux155),.in6(mux156),.in7(mux157),.in8(mux158),.in9(mux159),.in10(mux183),.in11(mux184),.in12(mux185),.in13(mux186),.in14(mux187),.in15(mux211),.in16(mux212),.in17(mux213),.in18(mux214),.in19(mux215),.in20(mux239),.in21(mux240),.in22(mux241),.in23(mux242),.in24(mux243), .bias(bias), .clk(clk), .out(muxin111));
 
Conv5D  Conv5D112(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux128),.in1(mux129),.in2(mux130),.in3(mux131),.in4(mux132),.in5(mux156),.in6(mux157),.in7(mux158),.in8(mux159),.in9(mux160),.in10(mux184),.in11(mux185),.in12(mux186),.in13(mux187),.in14(mux188),.in15(mux212),.in16(mux213),.in17(mux214),.in18(mux215),.in19(mux216),.in20(mux240),.in21(mux241),.in22(mux242),.in23(mux243),.in24(mux244), .bias(bias), .clk(clk), .out(muxin112));
 
Conv5D  Conv5D113(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux129),.in1(mux130),.in2(mux131),.in3(mux132),.in4(mux133),.in5(mux157),.in6(mux158),.in7(mux159),.in8(mux160),.in9(mux161),.in10(mux185),.in11(mux186),.in12(mux187),.in13(mux188),.in14(mux189),.in15(mux213),.in16(mux214),.in17(mux215),.in18(mux216),.in19(mux217),.in20(mux241),.in21(mux242),.in22(mux243),.in23(mux244),.in24(mux245), .bias(bias), .clk(clk), .out(muxin113));
 
Conv5D  Conv5D114(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux130),.in1(mux131),.in2(mux132),.in3(mux133),.in4(mux134),.in5(mux158),.in6(mux159),.in7(mux160),.in8(mux161),.in9(mux162),.in10(mux186),.in11(mux187),.in12(mux188),.in13(mux189),.in14(mux190),.in15(mux214),.in16(mux215),.in17(mux216),.in18(mux217),.in19(mux218),.in20(mux242),.in21(mux243),.in22(mux244),.in23(mux245),.in24(mux246), .bias(bias), .clk(clk), .out(muxin114));
 
Conv5D  Conv5D115(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux131),.in1(mux132),.in2(mux133),.in3(mux134),.in4(mux135),.in5(mux159),.in6(mux160),.in7(mux161),.in8(mux162),.in9(mux163),.in10(mux187),.in11(mux188),.in12(mux189),.in13(mux190),.in14(mux191),.in15(mux215),.in16(mux216),.in17(mux217),.in18(mux218),.in19(mux219),.in20(mux243),.in21(mux244),.in22(mux245),.in23(mux246),.in24(mux247), .bias(bias), .clk(clk), .out(muxin115));
 
Conv5D  Conv5D116(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux132),.in1(mux133),.in2(mux134),.in3(mux135),.in4(mux136),.in5(mux160),.in6(mux161),.in7(mux162),.in8(mux163),.in9(mux164),.in10(mux188),.in11(mux189),.in12(mux190),.in13(mux191),.in14(mux192),.in15(mux216),.in16(mux217),.in17(mux218),.in18(mux219),.in19(mux220),.in20(mux244),.in21(mux245),.in22(mux246),.in23(mux247),.in24(mux248), .bias(bias), .clk(clk), .out(muxin116));
 
Conv5D  Conv5D117(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux133),.in1(mux134),.in2(mux135),.in3(mux136),.in4(mux137),.in5(mux161),.in6(mux162),.in7(mux163),.in8(mux164),.in9(mux165),.in10(mux189),.in11(mux190),.in12(mux191),.in13(mux192),.in14(mux193),.in15(mux217),.in16(mux218),.in17(mux219),.in18(mux220),.in19(mux221),.in20(mux245),.in21(mux246),.in22(mux247),.in23(mux248),.in24(mux249), .bias(bias), .clk(clk), .out(muxin117));
 
Conv5D  Conv5D118(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux134),.in1(mux135),.in2(mux136),.in3(mux137),.in4(mux138),.in5(mux162),.in6(mux163),.in7(mux164),.in8(mux165),.in9(mux166),.in10(mux190),.in11(mux191),.in12(mux192),.in13(mux193),.in14(mux194),.in15(mux218),.in16(mux219),.in17(mux220),.in18(mux221),.in19(mux222),.in20(mux246),.in21(mux247),.in22(mux248),.in23(mux249),.in24(mux250), .bias(bias), .clk(clk), .out(muxin118));
 
Conv5D  Conv5D119(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux135),.in1(mux136),.in2(mux137),.in3(mux138),.in4(mux139),.in5(mux163),.in6(mux164),.in7(mux165),.in8(mux166),.in9(mux167),.in10(mux191),.in11(mux192),.in12(mux193),.in13(mux194),.in14(mux195),.in15(mux219),.in16(mux220),.in17(mux221),.in18(mux222),.in19(mux223),.in20(mux247),.in21(mux248),.in22(mux249),.in23(mux250),.in24(mux251), .bias(bias), .clk(clk), .out(muxin119));
 
Conv5D  Conv5D120(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux140),.in1(mux141),.in2(mux142),.in3(mux143),.in4(mux144),.in5(mux168),.in6(mux169),.in7(mux170),.in8(mux171),.in9(mux172),.in10(mux196),.in11(mux197),.in12(mux198),.in13(mux199),.in14(mux200),.in15(mux224),.in16(mux225),.in17(mux226),.in18(mux227),.in19(mux228),.in20(mux252),.in21(mux253),.in22(mux254),.in23(mux255),.in24(mux256), .bias(bias), .clk(clk), .out(muxin120));
 
Conv5D  Conv5D121(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux141),.in1(mux142),.in2(mux143),.in3(mux144),.in4(mux145),.in5(mux169),.in6(mux170),.in7(mux171),.in8(mux172),.in9(mux173),.in10(mux197),.in11(mux198),.in12(mux199),.in13(mux200),.in14(mux201),.in15(mux225),.in16(mux226),.in17(mux227),.in18(mux228),.in19(mux229),.in20(mux253),.in21(mux254),.in22(mux255),.in23(mux256),.in24(mux257), .bias(bias), .clk(clk), .out(muxin121));
 
Conv5D  Conv5D122(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux142),.in1(mux143),.in2(mux144),.in3(mux145),.in4(mux146),.in5(mux170),.in6(mux171),.in7(mux172),.in8(mux173),.in9(mux174),.in10(mux198),.in11(mux199),.in12(mux200),.in13(mux201),.in14(mux202),.in15(mux226),.in16(mux227),.in17(mux228),.in18(mux229),.in19(mux230),.in20(mux254),.in21(mux255),.in22(mux256),.in23(mux257),.in24(mux258), .bias(bias), .clk(clk), .out(muxin122));
 
Conv5D  Conv5D123(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux143),.in1(mux144),.in2(mux145),.in3(mux146),.in4(mux147),.in5(mux171),.in6(mux172),.in7(mux173),.in8(mux174),.in9(mux175),.in10(mux199),.in11(mux200),.in12(mux201),.in13(mux202),.in14(mux203),.in15(mux227),.in16(mux228),.in17(mux229),.in18(mux230),.in19(mux231),.in20(mux255),.in21(mux256),.in22(mux257),.in23(mux258),.in24(mux259), .bias(bias), .clk(clk), .out(muxin123));
 
Conv5D  Conv5D124(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux144),.in1(mux145),.in2(mux146),.in3(mux147),.in4(mux148),.in5(mux172),.in6(mux173),.in7(mux174),.in8(mux175),.in9(mux176),.in10(mux200),.in11(mux201),.in12(mux202),.in13(mux203),.in14(mux204),.in15(mux228),.in16(mux229),.in17(mux230),.in18(mux231),.in19(mux232),.in20(mux256),.in21(mux257),.in22(mux258),.in23(mux259),.in24(mux260), .bias(bias), .clk(clk), .out(muxin124));
 
Conv5D  Conv5D125(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux145),.in1(mux146),.in2(mux147),.in3(mux148),.in4(mux149),.in5(mux173),.in6(mux174),.in7(mux175),.in8(mux176),.in9(mux177),.in10(mux201),.in11(mux202),.in12(mux203),.in13(mux204),.in14(mux205),.in15(mux229),.in16(mux230),.in17(mux231),.in18(mux232),.in19(mux233),.in20(mux257),.in21(mux258),.in22(mux259),.in23(mux260),.in24(mux261), .bias(bias), .clk(clk), .out(muxin125));
 
Conv5D  Conv5D126(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux146),.in1(mux147),.in2(mux148),.in3(mux149),.in4(mux150),.in5(mux174),.in6(mux175),.in7(mux176),.in8(mux177),.in9(mux178),.in10(mux202),.in11(mux203),.in12(mux204),.in13(mux205),.in14(mux206),.in15(mux230),.in16(mux231),.in17(mux232),.in18(mux233),.in19(mux234),.in20(mux258),.in21(mux259),.in22(mux260),.in23(mux261),.in24(mux262), .bias(bias), .clk(clk), .out(muxin126));
 
Conv5D  Conv5D127(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux147),.in1(mux148),.in2(mux149),.in3(mux150),.in4(mux151),.in5(mux175),.in6(mux176),.in7(mux177),.in8(mux178),.in9(mux179),.in10(mux203),.in11(mux204),.in12(mux205),.in13(mux206),.in14(mux207),.in15(mux231),.in16(mux232),.in17(mux233),.in18(mux234),.in19(mux235),.in20(mux259),.in21(mux260),.in22(mux261),.in23(mux262),.in24(mux263), .bias(bias), .clk(clk), .out(muxin127));
 
Conv5D  Conv5D128(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux148),.in1(mux149),.in2(mux150),.in3(mux151),.in4(mux152),.in5(mux176),.in6(mux177),.in7(mux178),.in8(mux179),.in9(mux180),.in10(mux204),.in11(mux205),.in12(mux206),.in13(mux207),.in14(mux208),.in15(mux232),.in16(mux233),.in17(mux234),.in18(mux235),.in19(mux236),.in20(mux260),.in21(mux261),.in22(mux262),.in23(mux263),.in24(mux264), .bias(bias), .clk(clk), .out(muxin128));
 
Conv5D  Conv5D129(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux149),.in1(mux150),.in2(mux151),.in3(mux152),.in4(mux153),.in5(mux177),.in6(mux178),.in7(mux179),.in8(mux180),.in9(mux181),.in10(mux205),.in11(mux206),.in12(mux207),.in13(mux208),.in14(mux209),.in15(mux233),.in16(mux234),.in17(mux235),.in18(mux236),.in19(mux237),.in20(mux261),.in21(mux262),.in22(mux263),.in23(mux264),.in24(mux265), .bias(bias), .clk(clk), .out(muxin129));
 
Conv5D  Conv5D130(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux150),.in1(mux151),.in2(mux152),.in3(mux153),.in4(mux154),.in5(mux178),.in6(mux179),.in7(mux180),.in8(mux181),.in9(mux182),.in10(mux206),.in11(mux207),.in12(mux208),.in13(mux209),.in14(mux210),.in15(mux234),.in16(mux235),.in17(mux236),.in18(mux237),.in19(mux238),.in20(mux262),.in21(mux263),.in22(mux264),.in23(mux265),.in24(mux266), .bias(bias), .clk(clk), .out(muxin130));
 
Conv5D  Conv5D131(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux151),.in1(mux152),.in2(mux153),.in3(mux154),.in4(mux155),.in5(mux179),.in6(mux180),.in7(mux181),.in8(mux182),.in9(mux183),.in10(mux207),.in11(mux208),.in12(mux209),.in13(mux210),.in14(mux211),.in15(mux235),.in16(mux236),.in17(mux237),.in18(mux238),.in19(mux239),.in20(mux263),.in21(mux264),.in22(mux265),.in23(mux266),.in24(mux267), .bias(bias), .clk(clk), .out(muxin131));
 
Conv5D  Conv5D132(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux152),.in1(mux153),.in2(mux154),.in3(mux155),.in4(mux156),.in5(mux180),.in6(mux181),.in7(mux182),.in8(mux183),.in9(mux184),.in10(mux208),.in11(mux209),.in12(mux210),.in13(mux211),.in14(mux212),.in15(mux236),.in16(mux237),.in17(mux238),.in18(mux239),.in19(mux240),.in20(mux264),.in21(mux265),.in22(mux266),.in23(mux267),.in24(mux268), .bias(bias), .clk(clk), .out(muxin132));
 
Conv5D  Conv5D133(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux153),.in1(mux154),.in2(mux155),.in3(mux156),.in4(mux157),.in5(mux181),.in6(mux182),.in7(mux183),.in8(mux184),.in9(mux185),.in10(mux209),.in11(mux210),.in12(mux211),.in13(mux212),.in14(mux213),.in15(mux237),.in16(mux238),.in17(mux239),.in18(mux240),.in19(mux241),.in20(mux265),.in21(mux266),.in22(mux267),.in23(mux268),.in24(mux269), .bias(bias), .clk(clk), .out(muxin133));
 
Conv5D  Conv5D134(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux154),.in1(mux155),.in2(mux156),.in3(mux157),.in4(mux158),.in5(mux182),.in6(mux183),.in7(mux184),.in8(mux185),.in9(mux186),.in10(mux210),.in11(mux211),.in12(mux212),.in13(mux213),.in14(mux214),.in15(mux238),.in16(mux239),.in17(mux240),.in18(mux241),.in19(mux242),.in20(mux266),.in21(mux267),.in22(mux268),.in23(mux269),.in24(mux270), .bias(bias), .clk(clk), .out(muxin134));
 
Conv5D  Conv5D135(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux155),.in1(mux156),.in2(mux157),.in3(mux158),.in4(mux159),.in5(mux183),.in6(mux184),.in7(mux185),.in8(mux186),.in9(mux187),.in10(mux211),.in11(mux212),.in12(mux213),.in13(mux214),.in14(mux215),.in15(mux239),.in16(mux240),.in17(mux241),.in18(mux242),.in19(mux243),.in20(mux267),.in21(mux268),.in22(mux269),.in23(mux270),.in24(mux271), .bias(bias), .clk(clk), .out(muxin135));
 
Conv5D  Conv5D136(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux156),.in1(mux157),.in2(mux158),.in3(mux159),.in4(mux160),.in5(mux184),.in6(mux185),.in7(mux186),.in8(mux187),.in9(mux188),.in10(mux212),.in11(mux213),.in12(mux214),.in13(mux215),.in14(mux216),.in15(mux240),.in16(mux241),.in17(mux242),.in18(mux243),.in19(mux244),.in20(mux268),.in21(mux269),.in22(mux270),.in23(mux271),.in24(mux272), .bias(bias), .clk(clk), .out(muxin136));
 
Conv5D  Conv5D137(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux157),.in1(mux158),.in2(mux159),.in3(mux160),.in4(mux161),.in5(mux185),.in6(mux186),.in7(mux187),.in8(mux188),.in9(mux189),.in10(mux213),.in11(mux214),.in12(mux215),.in13(mux216),.in14(mux217),.in15(mux241),.in16(mux242),.in17(mux243),.in18(mux244),.in19(mux245),.in20(mux269),.in21(mux270),.in22(mux271),.in23(mux272),.in24(mux273), .bias(bias), .clk(clk), .out(muxin137));
 
Conv5D  Conv5D138(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux158),.in1(mux159),.in2(mux160),.in3(mux161),.in4(mux162),.in5(mux186),.in6(mux187),.in7(mux188),.in8(mux189),.in9(mux190),.in10(mux214),.in11(mux215),.in12(mux216),.in13(mux217),.in14(mux218),.in15(mux242),.in16(mux243),.in17(mux244),.in18(mux245),.in19(mux246),.in20(mux270),.in21(mux271),.in22(mux272),.in23(mux273),.in24(mux274), .bias(bias), .clk(clk), .out(muxin138));
 
Conv5D  Conv5D139(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux159),.in1(mux160),.in2(mux161),.in3(mux162),.in4(mux163),.in5(mux187),.in6(mux188),.in7(mux189),.in8(mux190),.in9(mux191),.in10(mux215),.in11(mux216),.in12(mux217),.in13(mux218),.in14(mux219),.in15(mux243),.in16(mux244),.in17(mux245),.in18(mux246),.in19(mux247),.in20(mux271),.in21(mux272),.in22(mux273),.in23(mux274),.in24(mux275), .bias(bias), .clk(clk), .out(muxin139));
 
Conv5D  Conv5D140(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux160),.in1(mux161),.in2(mux162),.in3(mux163),.in4(mux164),.in5(mux188),.in6(mux189),.in7(mux190),.in8(mux191),.in9(mux192),.in10(mux216),.in11(mux217),.in12(mux218),.in13(mux219),.in14(mux220),.in15(mux244),.in16(mux245),.in17(mux246),.in18(mux247),.in19(mux248),.in20(mux272),.in21(mux273),.in22(mux274),.in23(mux275),.in24(mux276), .bias(bias), .clk(clk), .out(muxin140));
 
Conv5D  Conv5D141(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux161),.in1(mux162),.in2(mux163),.in3(mux164),.in4(mux165),.in5(mux189),.in6(mux190),.in7(mux191),.in8(mux192),.in9(mux193),.in10(mux217),.in11(mux218),.in12(mux219),.in13(mux220),.in14(mux221),.in15(mux245),.in16(mux246),.in17(mux247),.in18(mux248),.in19(mux249),.in20(mux273),.in21(mux274),.in22(mux275),.in23(mux276),.in24(mux277), .bias(bias), .clk(clk), .out(muxin141));
 
Conv5D  Conv5D142(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux162),.in1(mux163),.in2(mux164),.in3(mux165),.in4(mux166),.in5(mux190),.in6(mux191),.in7(mux192),.in8(mux193),.in9(mux194),.in10(mux218),.in11(mux219),.in12(mux220),.in13(mux221),.in14(mux222),.in15(mux246),.in16(mux247),.in17(mux248),.in18(mux249),.in19(mux250),.in20(mux274),.in21(mux275),.in22(mux276),.in23(mux277),.in24(mux278), .bias(bias), .clk(clk), .out(muxin142));
 
Conv5D  Conv5D143(.weight0(weight0),.weight1(weight1),.weight2(weight2),.weight3(weight3),.weight4(weight4),.weight5(weight5),.weight6(weight6),.weight7(weight7),.weight8(weight8),.weight9(weight9),.weight10(weight10),.weight11(weight11),.weight12(weight12),.weight13(weight13),.weight14(weight14),.weight15(weight15),.weight16(weight16),.weight17(weight17),.weight18(weight18),.weight19(weight19),.weight20(weight20),.weight21(weight21),.weight22(weight22),.weight23(weight23),.weight24(weight24),.in0(mux163),.in1(mux164),.in2(mux165),.in3(mux166),.in4(mux167),.in5(mux191),.in6(mux192),.in7(mux193),.in8(mux194),.in9(mux195),.in10(mux219),.in11(mux220),.in12(mux221),.in13(mux222),.in14(mux223),.in15(mux247),.in16(mux248),.in17(mux249),.in18(mux250),.in19(mux251),.in20(mux275),.in21(mux276),.in22(mux277),.in23(mux278),.in24(mux279), .bias(bias), .clk(clk), .out(muxin143));
 



endmodule

module mux42(a,b,c,d,sel,out);

input [7:0] a;
input [7:0] b;
input [7:0] c;
input [7:0] d;
input [1:0] sel;
output [7:0] out;
reg [7:0] out;

always @(*)
begin
	case(sel)
		2'b00:
			out = a;
		2'b01:
			out = b;
		2'b10:
			out = c;
		2'b11:
			out = d;
	endcase
end

endmodule

module demux42(a,b,c,d,sel,out);

output [7:0] a;
output [7:0] b;
output [7:0] c;
output [7:0] d;
reg [7:0] a;
reg [7:0] b;
reg [7:0] c;
reg [7:0] d;
input [1:0] sel;
input [7:0] out;

always @(*)
begin
	case(sel)
		2'b00:
			a <= out;
		2'b01:
			b <= out;
		2'b10:
			c <= out;
		2'b11:
			d <= out;
	endcase
end
endmodule