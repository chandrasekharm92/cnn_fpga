`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    20:58:17 11/02/2017 
// Design Name: 
// Module Name:    testbench 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module testbench();
reg [7:0]weight[24:0];
reg [7:0]weight2l[143:0];
reg [7:0]in[783:0];
reg [7:0]bias;
wire [7:0] out;
reg start;
reg clk;
wire ready;
wire [7:0]conv[575:0];

integer i;
initial begin
	start = 0;
	for(i=0;i<25;i=i+1)begin
		weight[i] = 8'd1;
	end
	for(i=0;i<144;i=i+1)begin
		weight2l[i] = 8'd1;
	end
	for(i=0;i<784;i=i+1)begin
		in[i] = i;
	end
	bias = 8'b1;
	clk = 1'b0;
	#10 start = 1;
	#15 start = 0;	
end

cnn cnn1(
 .weight1l0(weight[0]),.weight1l1(weight[1]),.weight1l2(weight[2]),.weight1l3(weight[3]),.weight1l4(weight[4]),.weight1l5(weight[5]),.weight1l6(weight[6]),.weight1l7(weight[7]),.weight1l8(weight[8]),.weight1l9(weight[9]),.weight1l10(weight[10]),.weight1l11(weight[11]),.weight1l12(weight[12]),.weight1l13(weight[13]),.weight1l14(weight[14]),.weight1l15(weight[15]),.weight1l16(weight[16]),.weight1l17(weight[17]),.weight1l18(weight[18]),.weight1l19(weight[19]),.weight1l20(weight[20]),.weight1l21(weight[21]),.weight1l22(weight[22]),.weight1l23(weight[23]),.weight1l24(weight[24]),
.weight2l0(weight2l[0]),.weight2l1(weight2l[1]),.weight2l2(weight2l[2]),.weight2l3(weight2l[3]),.weight2l4(weight2l[4]),.weight2l5(weight2l[5]),.weight2l6(weight2l[6]),.weight2l7(weight2l[7]),.weight2l8(weight2l[8]),.weight2l9(weight2l[9]),.weight2l10(weight2l[10]),.weight2l11(weight2l[11]),.weight2l12(weight2l[12]),.weight2l13(weight2l[13]),.weight2l14(weight2l[14]),.weight2l15(weight2l[15]),.weight2l16(weight2l[16]),.weight2l17(weight2l[17]),.weight2l18(weight2l[18]),.weight2l19(weight2l[19]),.weight2l20(weight2l[20]),.weight2l21(weight2l[21]),.weight2l22(weight2l[22]),.weight2l23(weight2l[23]),.weight2l24(weight2l[24]),.weight2l25(weight2l[25]),.weight2l26(weight2l[26]),.weight2l27(weight2l[27]),.weight2l28(weight2l[28]),.weight2l29(weight2l[29]),.weight2l30(weight2l[30]),.weight2l31(weight2l[31]),.weight2l32(weight2l[32]),.weight2l33(weight2l[33]),.weight2l34(weight2l[34]),.weight2l35(weight2l[35]),.weight2l36(weight2l[36]),.weight2l37(weight2l[37]),.weight2l38(weight2l[38]),.weight2l39(weight2l[39]),.weight2l40(weight2l[40]),.weight2l41(weight2l[41]),.weight2l42(weight2l[42]),.weight2l43(weight2l[43]),.weight2l44(weight2l[44]),.weight2l45(weight2l[45]),.weight2l46(weight2l[46]),.weight2l47(weight2l[47]),.weight2l48(weight2l[48]),.weight2l49(weight2l[49]),.weight2l50(weight2l[50]),.weight2l51(weight2l[51]),.weight2l52(weight2l[52]),.weight2l53(weight2l[53]),.weight2l54(weight2l[54]),.weight2l55(weight2l[55]),.weight2l56(weight2l[56]),.weight2l57(weight2l[57]),.weight2l58(weight2l[58]),.weight2l59(weight2l[59]),.weight2l60(weight2l[60]),.weight2l61(weight2l[61]),.weight2l62(weight2l[62]),.weight2l63(weight2l[63]),.weight2l64(weight2l[64]),.weight2l65(weight2l[65]),.weight2l66(weight2l[66]),.weight2l67(weight2l[67]),.weight2l68(weight2l[68]),.weight2l69(weight2l[69]),.weight2l70(weight2l[70]),.weight2l71(weight2l[71]),.weight2l72(weight2l[72]),.weight2l73(weight2l[73]),.weight2l74(weight2l[74]),.weight2l75(weight2l[75]),.weight2l76(weight2l[76]),.weight2l77(weight2l[77]),.weight2l78(weight2l[78]),.weight2l79(weight2l[79]),.weight2l80(weight2l[80]),.weight2l81(weight2l[81]),.weight2l82(weight2l[82]),.weight2l83(weight2l[83]),.weight2l84(weight2l[84]),.weight2l85(weight2l[85]),.weight2l86(weight2l[86]),.weight2l87(weight2l[87]),.weight2l88(weight2l[88]),.weight2l89(weight2l[89]),.weight2l90(weight2l[90]),.weight2l91(weight2l[91]),.weight2l92(weight2l[92]),.weight2l93(weight2l[93]),.weight2l94(weight2l[94]),.weight2l95(weight2l[95]),.weight2l96(weight2l[96]),.weight2l97(weight2l[97]),.weight2l98(weight2l[98]),.weight2l99(weight2l[99]),.weight2l100(weight2l[100]),.weight2l101(weight2l[101]),.weight2l102(weight2l[102]),.weight2l103(weight2l[103]),.weight2l104(weight2l[104]),.weight2l105(weight2l[105]),.weight2l106(weight2l[106]),.weight2l107(weight2l[107]),.weight2l108(weight2l[108]),.weight2l109(weight2l[109]),.weight2l110(weight2l[110]),.weight2l111(weight2l[111]),.weight2l112(weight2l[112]),.weight2l113(weight2l[113]),.weight2l114(weight2l[114]),.weight2l115(weight2l[115]),.weight2l116(weight2l[116]),.weight2l117(weight2l[117]),.weight2l118(weight2l[118]),.weight2l119(weight2l[119]),.weight2l120(weight2l[120]),.weight2l121(weight2l[121]),.weight2l122(weight2l[122]),.weight2l123(weight2l[123]),.weight2l124(weight2l[124]),.weight2l125(weight2l[125]),.weight2l126(weight2l[126]),.weight2l127(weight2l[127]),.weight2l128(weight2l[128]),.weight2l129(weight2l[129]),.weight2l130(weight2l[130]),.weight2l131(weight2l[131]),.weight2l132(weight2l[132]),.weight2l133(weight2l[133]),.weight2l134(weight2l[134]),.weight2l135(weight2l[135]),.weight2l136(weight2l[136]),.weight2l137(weight2l[137]),.weight2l138(weight2l[138]),.weight2l139(weight2l[139]),.weight2l140(weight2l[140]),.weight2l141(weight2l[141]),.weight2l142(weight2l[142]),.weight2l143(weight2l[143]),
 .in0(in[0]),.in1(in[1]),.in2(in[2]),.in3(in[3]),.in4(in[4]),.in5(in[5]),.in6(in[6]),.in7(in[7]),.in8(in[8]),.in9(in[9]),.in10(in[10]),.in11(in[11]),.in12(in[12]),.in13(in[13]),.in14(in[14]),.in15(in[15]),.in16(in[16]),.in17(in[17]),.in18(in[18]),.in19(in[19]),.in20(in[20]),.in21(in[21]),.in22(in[22]),.in23(in[23]),.in24(in[24]),.in25(in[25]),.in26(in[26]),.in27(in[27]),.in28(in[28]),.in29(in[29]),.in30(in[30]),.in31(in[31]),.in32(in[32]),.in33(in[33]),.in34(in[34]),.in35(in[35]),.in36(in[36]),.in37(in[37]),.in38(in[38]),.in39(in[39]),.in40(in[40]),.in41(in[41]),.in42(in[42]),.in43(in[43]),.in44(in[44]),.in45(in[45]),.in46(in[46]),.in47(in[47]),.in48(in[48]),.in49(in[49]),.in50(in[50]),.in51(in[51]),.in52(in[52]),.in53(in[53]),.in54(in[54]),.in55(in[55]),.in56(in[56]),.in57(in[57]),.in58(in[58]),.in59(in[59]),.in60(in[60]),.in61(in[61]),.in62(in[62]),.in63(in[63]),.in64(in[64]),.in65(in[65]),.in66(in[66]),.in67(in[67]),.in68(in[68]),.in69(in[69]),.in70(in[70]),.in71(in[71]),.in72(in[72]),.in73(in[73]),.in74(in[74]),.in75(in[75]),.in76(in[76]),.in77(in[77]),.in78(in[78]),.in79(in[79]),.in80(in[80]),.in81(in[81]),.in82(in[82]),.in83(in[83]),.in84(in[84]),.in85(in[85]),.in86(in[86]),.in87(in[87]),.in88(in[88]),.in89(in[89]),.in90(in[90]),.in91(in[91]),.in92(in[92]),.in93(in[93]),.in94(in[94]),.in95(in[95]),.in96(in[96]),.in97(in[97]),.in98(in[98]),.in99(in[99]),.in100(in[100]),.in101(in[101]),.in102(in[102]),.in103(in[103]),.in104(in[104]),.in105(in[105]),.in106(in[106]),.in107(in[107]),.in108(in[108]),.in109(in[109]),.in110(in[110]),.in111(in[111]),.in112(in[112]),.in113(in[113]),.in114(in[114]),.in115(in[115]),.in116(in[116]),.in117(in[117]),.in118(in[118]),.in119(in[119]),.in120(in[120]),.in121(in[121]),.in122(in[122]),.in123(in[123]),.in124(in[124]),.in125(in[125]),.in126(in[126]),.in127(in[127]),.in128(in[128]),.in129(in[129]),.in130(in[130]),.in131(in[131]),.in132(in[132]),.in133(in[133]),.in134(in[134]),.in135(in[135]),.in136(in[136]),.in137(in[137]),.in138(in[138]),.in139(in[139]),.in140(in[140]),.in141(in[141]),.in142(in[142]),.in143(in[143]),.in144(in[144]),.in145(in[145]),.in146(in[146]),.in147(in[147]),.in148(in[148]),.in149(in[149]),.in150(in[150]),.in151(in[151]),.in152(in[152]),.in153(in[153]),.in154(in[154]),.in155(in[155]),.in156(in[156]),.in157(in[157]),.in158(in[158]),.in159(in[159]),.in160(in[160]),.in161(in[161]),.in162(in[162]),.in163(in[163]),.in164(in[164]),.in165(in[165]),.in166(in[166]),.in167(in[167]),.in168(in[168]),.in169(in[169]),.in170(in[170]),.in171(in[171]),.in172(in[172]),.in173(in[173]),.in174(in[174]),.in175(in[175]),.in176(in[176]),.in177(in[177]),.in178(in[178]),.in179(in[179]),.in180(in[180]),.in181(in[181]),.in182(in[182]),.in183(in[183]),.in184(in[184]),.in185(in[185]),.in186(in[186]),.in187(in[187]),.in188(in[188]),.in189(in[189]),.in190(in[190]),.in191(in[191]),.in192(in[192]),.in193(in[193]),.in194(in[194]),.in195(in[195]),.in196(in[196]),.in197(in[197]),.in198(in[198]),.in199(in[199]),.in200(in[200]),.in201(in[201]),.in202(in[202]),.in203(in[203]),.in204(in[204]),.in205(in[205]),.in206(in[206]),.in207(in[207]),.in208(in[208]),.in209(in[209]),.in210(in[210]),.in211(in[211]),.in212(in[212]),.in213(in[213]),.in214(in[214]),.in215(in[215]),.in216(in[216]),.in217(in[217]),.in218(in[218]),.in219(in[219]),.in220(in[220]),.in221(in[221]),.in222(in[222]),.in223(in[223]),.in224(in[224]),.in225(in[225]),.in226(in[226]),.in227(in[227]),.in228(in[228]),.in229(in[229]),.in230(in[230]),.in231(in[231]),.in232(in[232]),.in233(in[233]),.in234(in[234]),.in235(in[235]),.in236(in[236]),.in237(in[237]),.in238(in[238]),.in239(in[239]),.in240(in[240]),.in241(in[241]),.in242(in[242]),.in243(in[243]),.in244(in[244]),.in245(in[245]),.in246(in[246]),.in247(in[247]),.in248(in[248]),.in249(in[249]),.in250(in[250]),.in251(in[251]),.in252(in[252]),.in253(in[253]),.in254(in[254]),.in255(in[255]),.in256(in[256]),.in257(in[257]),.in258(in[258]),.in259(in[259]),.in260(in[260]),.in261(in[261]),.in262(in[262]),.in263(in[263]),.in264(in[264]),.in265(in[265]),.in266(in[266]),.in267(in[267]),.in268(in[268]),.in269(in[269]),.in270(in[270]),.in271(in[271]),.in272(in[272]),.in273(in[273]),.in274(in[274]),.in275(in[275]),.in276(in[276]),.in277(in[277]),.in278(in[278]),.in279(in[279]),.in280(in[280]),.in281(in[281]),.in282(in[282]),.in283(in[283]),.in284(in[284]),.in285(in[285]),.in286(in[286]),.in287(in[287]),.in288(in[288]),.in289(in[289]),.in290(in[290]),.in291(in[291]),.in292(in[292]),.in293(in[293]),.in294(in[294]),.in295(in[295]),.in296(in[296]),.in297(in[297]),.in298(in[298]),.in299(in[299]),.in300(in[300]),.in301(in[301]),.in302(in[302]),.in303(in[303]),.in304(in[304]),.in305(in[305]),.in306(in[306]),.in307(in[307]),.in308(in[308]),.in309(in[309]),.in310(in[310]),.in311(in[311]),.in312(in[312]),.in313(in[313]),.in314(in[314]),.in315(in[315]),.in316(in[316]),.in317(in[317]),.in318(in[318]),.in319(in[319]),.in320(in[320]),.in321(in[321]),.in322(in[322]),.in323(in[323]),.in324(in[324]),.in325(in[325]),.in326(in[326]),.in327(in[327]),.in328(in[328]),.in329(in[329]),.in330(in[330]),.in331(in[331]),.in332(in[332]),.in333(in[333]),.in334(in[334]),.in335(in[335]),.in336(in[336]),.in337(in[337]),.in338(in[338]),.in339(in[339]),.in340(in[340]),.in341(in[341]),.in342(in[342]),.in343(in[343]),.in344(in[344]),.in345(in[345]),.in346(in[346]),.in347(in[347]),.in348(in[348]),.in349(in[349]),.in350(in[350]),.in351(in[351]),.in352(in[352]),.in353(in[353]),.in354(in[354]),.in355(in[355]),.in356(in[356]),.in357(in[357]),.in358(in[358]),.in359(in[359]),.in360(in[360]),.in361(in[361]),.in362(in[362]),.in363(in[363]),.in364(in[364]),.in365(in[365]),.in366(in[366]),.in367(in[367]),.in368(in[368]),.in369(in[369]),.in370(in[370]),.in371(in[371]),.in372(in[372]),.in373(in[373]),.in374(in[374]),.in375(in[375]),.in376(in[376]),.in377(in[377]),.in378(in[378]),.in379(in[379]),.in380(in[380]),.in381(in[381]),.in382(in[382]),.in383(in[383]),.in384(in[384]),.in385(in[385]),.in386(in[386]),.in387(in[387]),.in388(in[388]),.in389(in[389]),.in390(in[390]),.in391(in[391]),.in392(in[392]),.in393(in[393]),.in394(in[394]),.in395(in[395]),.in396(in[396]),.in397(in[397]),.in398(in[398]),.in399(in[399]),.in400(in[400]),.in401(in[401]),.in402(in[402]),.in403(in[403]),.in404(in[404]),.in405(in[405]),.in406(in[406]),.in407(in[407]),.in408(in[408]),.in409(in[409]),.in410(in[410]),.in411(in[411]),.in412(in[412]),.in413(in[413]),.in414(in[414]),.in415(in[415]),.in416(in[416]),.in417(in[417]),.in418(in[418]),.in419(in[419]),.in420(in[420]),.in421(in[421]),.in422(in[422]),.in423(in[423]),.in424(in[424]),.in425(in[425]),.in426(in[426]),.in427(in[427]),.in428(in[428]),.in429(in[429]),.in430(in[430]),.in431(in[431]),.in432(in[432]),.in433(in[433]),.in434(in[434]),.in435(in[435]),.in436(in[436]),.in437(in[437]),.in438(in[438]),.in439(in[439]),.in440(in[440]),.in441(in[441]),.in442(in[442]),.in443(in[443]),.in444(in[444]),.in445(in[445]),.in446(in[446]),.in447(in[447]),.in448(in[448]),.in449(in[449]),.in450(in[450]),.in451(in[451]),.in452(in[452]),.in453(in[453]),.in454(in[454]),.in455(in[455]),.in456(in[456]),.in457(in[457]),.in458(in[458]),.in459(in[459]),.in460(in[460]),.in461(in[461]),.in462(in[462]),.in463(in[463]),.in464(in[464]),.in465(in[465]),.in466(in[466]),.in467(in[467]),.in468(in[468]),.in469(in[469]),.in470(in[470]),.in471(in[471]),.in472(in[472]),.in473(in[473]),.in474(in[474]),.in475(in[475]),.in476(in[476]),.in477(in[477]),.in478(in[478]),.in479(in[479]),.in480(in[480]),.in481(in[481]),.in482(in[482]),.in483(in[483]),.in484(in[484]),.in485(in[485]),.in486(in[486]),.in487(in[487]),.in488(in[488]),.in489(in[489]),.in490(in[490]),.in491(in[491]),.in492(in[492]),.in493(in[493]),.in494(in[494]),.in495(in[495]),.in496(in[496]),.in497(in[497]),.in498(in[498]),.in499(in[499]),.in500(in[500]),.in501(in[501]),.in502(in[502]),.in503(in[503]),.in504(in[504]),.in505(in[505]),.in506(in[506]),.in507(in[507]),.in508(in[508]),.in509(in[509]),.in510(in[510]),.in511(in[511]),.in512(in[512]),.in513(in[513]),.in514(in[514]),.in515(in[515]),.in516(in[516]),.in517(in[517]),.in518(in[518]),.in519(in[519]),.in520(in[520]),.in521(in[521]),.in522(in[522]),.in523(in[523]),.in524(in[524]),.in525(in[525]),.in526(in[526]),.in527(in[527]),.in528(in[528]),.in529(in[529]),.in530(in[530]),.in531(in[531]),.in532(in[532]),.in533(in[533]),.in534(in[534]),.in535(in[535]),.in536(in[536]),.in537(in[537]),.in538(in[538]),.in539(in[539]),.in540(in[540]),.in541(in[541]),.in542(in[542]),.in543(in[543]),.in544(in[544]),.in545(in[545]),.in546(in[546]),.in547(in[547]),.in548(in[548]),.in549(in[549]),.in550(in[550]),.in551(in[551]),.in552(in[552]),.in553(in[553]),.in554(in[554]),.in555(in[555]),.in556(in[556]),.in557(in[557]),.in558(in[558]),.in559(in[559]),.in560(in[560]),.in561(in[561]),.in562(in[562]),.in563(in[563]),.in564(in[564]),.in565(in[565]),.in566(in[566]),.in567(in[567]),.in568(in[568]),.in569(in[569]),.in570(in[570]),.in571(in[571]),.in572(in[572]),.in573(in[573]),.in574(in[574]),.in575(in[575]),.in576(in[576]),.in577(in[577]),.in578(in[578]),.in579(in[579]),.in580(in[580]),.in581(in[581]),.in582(in[582]),.in583(in[583]),.in584(in[584]),.in585(in[585]),.in586(in[586]),.in587(in[587]),.in588(in[588]),.in589(in[589]),.in590(in[590]),.in591(in[591]),.in592(in[592]),.in593(in[593]),.in594(in[594]),.in595(in[595]),.in596(in[596]),.in597(in[597]),.in598(in[598]),.in599(in[599]),.in600(in[600]),.in601(in[601]),.in602(in[602]),.in603(in[603]),.in604(in[604]),.in605(in[605]),.in606(in[606]),.in607(in[607]),.in608(in[608]),.in609(in[609]),.in610(in[610]),.in611(in[611]),.in612(in[612]),.in613(in[613]),.in614(in[614]),.in615(in[615]),.in616(in[616]),.in617(in[617]),.in618(in[618]),.in619(in[619]),.in620(in[620]),.in621(in[621]),.in622(in[622]),.in623(in[623]),.in624(in[624]),.in625(in[625]),.in626(in[626]),.in627(in[627]),.in628(in[628]),.in629(in[629]),.in630(in[630]),.in631(in[631]),.in632(in[632]),.in633(in[633]),.in634(in[634]),.in635(in[635]),.in636(in[636]),.in637(in[637]),.in638(in[638]),.in639(in[639]),.in640(in[640]),.in641(in[641]),.in642(in[642]),.in643(in[643]),.in644(in[644]),.in645(in[645]),.in646(in[646]),.in647(in[647]),.in648(in[648]),.in649(in[649]),.in650(in[650]),.in651(in[651]),.in652(in[652]),.in653(in[653]),.in654(in[654]),.in655(in[655]),.in656(in[656]),.in657(in[657]),.in658(in[658]),.in659(in[659]),.in660(in[660]),.in661(in[661]),.in662(in[662]),.in663(in[663]),.in664(in[664]),.in665(in[665]),.in666(in[666]),.in667(in[667]),.in668(in[668]),.in669(in[669]),.in670(in[670]),.in671(in[671]),.in672(in[672]),.in673(in[673]),.in674(in[674]),.in675(in[675]),.in676(in[676]),.in677(in[677]),.in678(in[678]),.in679(in[679]),.in680(in[680]),.in681(in[681]),.in682(in[682]),.in683(in[683]),.in684(in[684]),.in685(in[685]),.in686(in[686]),.in687(in[687]),.in688(in[688]),.in689(in[689]),.in690(in[690]),.in691(in[691]),.in692(in[692]),.in693(in[693]),.in694(in[694]),.in695(in[695]),.in696(in[696]),.in697(in[697]),.in698(in[698]),.in699(in[699]),.in700(in[700]),.in701(in[701]),.in702(in[702]),.in703(in[703]),.in704(in[704]),.in705(in[705]),.in706(in[706]),.in707(in[707]),.in708(in[708]),.in709(in[709]),.in710(in[710]),.in711(in[711]),.in712(in[712]),.in713(in[713]),.in714(in[714]),.in715(in[715]),.in716(in[716]),.in717(in[717]),.in718(in[718]),.in719(in[719]),.in720(in[720]),.in721(in[721]),.in722(in[722]),.in723(in[723]),.in724(in[724]),.in725(in[725]),.in726(in[726]),.in727(in[727]),.in728(in[728]),.in729(in[729]),.in730(in[730]),.in731(in[731]),.in732(in[732]),.in733(in[733]),.in734(in[734]),.in735(in[735]),.in736(in[736]),.in737(in[737]),.in738(in[738]),.in739(in[739]),.in740(in[740]),.in741(in[741]),.in742(in[742]),.in743(in[743]),.in744(in[744]),.in745(in[745]),.in746(in[746]),.in747(in[747]),.in748(in[748]),.in749(in[749]),.in750(in[750]),.in751(in[751]),.in752(in[752]),.in753(in[753]),.in754(in[754]),.in755(in[755]),.in756(in[756]),.in757(in[757]),.in758(in[758]),.in759(in[759]),.in760(in[760]),.in761(in[761]),.in762(in[762]),.in763(in[763]),.in764(in[764]),.in765(in[765]),.in766(in[766]),.in767(in[767]),.in768(in[768]),.in769(in[769]),.in770(in[770]),.in771(in[771]),.in772(in[772]),.in773(in[773]),.in774(in[774]),.in775(in[775]),.in776(in[776]),.in777(in[777]),.in778(in[778]),.in779(in[779]),.in780(in[780]),.in781(in[781]),.in782(in[782]),.in783(in[783]),.clk(clk),.ready(ready),.start(start),.bias(bias),.out(out)
);

/*poolinglayer poolinglayer1(
.out0(conv[0]),.out1(conv[1]),.out2(conv[2]),.out3(conv[3]),.out4(conv[4]),.out5(conv[5]),.out6(conv[6]),.out7(conv[7]),.out8(conv[8]),.out9(conv[9]),.out10(conv[10]),.out11(conv[11]),.out12(conv[12]),.out13(conv[13]),.out14(conv[14]),.out15(conv[15]),.out16(conv[16]),.out17(conv[17]),.out18(conv[18]),.out19(conv[19]),.out20(conv[20]),.out21(conv[21]),.out22(conv[22]),.out23(conv[23]),.out24(conv[24]),.out25(conv[25]),.out26(conv[26]),.out27(conv[27]),.out28(conv[28]),.out29(conv[29]),.out30(conv[30]),.out31(conv[31]),.out32(conv[32]),.out33(conv[33]),.out34(conv[34]),.out35(conv[35]),.out36(conv[36]),.out37(conv[37]),.out38(conv[38]),.out39(conv[39]),.out40(conv[40]),.out41(conv[41]),.out42(conv[42]),.out43(conv[43]),.out44(conv[44]),.out45(conv[45]),.out46(conv[46]),.out47(conv[47]),.out48(conv[48]),.out49(conv[49]),.out50(conv[50]),.out51(conv[51]),.out52(conv[52]),.out53(conv[53]),.out54(conv[54]),.out55(conv[55]),.out56(conv[56]),.out57(conv[57]),.out58(conv[58]),.out59(conv[59]),.out60(conv[60]),.out61(conv[61]),.out62(conv[62]),.out63(conv[63]),.out64(conv[64]),.out65(conv[65]),.out66(conv[66]),.out67(conv[67]),.out68(conv[68]),.out69(conv[69]),.out70(conv[70]),.out71(conv[71]),.out72(conv[72]),.out73(conv[73]),.out74(conv[74]),.out75(conv[75]),.out76(conv[76]),.out77(conv[77]),.out78(conv[78]),.out79(conv[79]),.out80(conv[80]),.out81(conv[81]),.out82(conv[82]),.out83(conv[83]),.out84(conv[84]),.out85(conv[85]),.out86(conv[86]),.out87(conv[87]),.out88(conv[88]),.out89(conv[89]),.out90(conv[90]),.out91(conv[91]),.out92(conv[92]),.out93(conv[93]),.out94(conv[94]),.out95(conv[95]),.out96(conv[96]),.out97(conv[97]),.out98(conv[98]),.out99(conv[99]),.out100(conv[100]),.out101(conv[101]),.out102(conv[102]),.out103(conv[103]),.out104(conv[104]),.out105(conv[105]),.out106(conv[106]),.out107(conv[107]),.out108(conv[108]),.out109(conv[109]),.out110(conv[110]),.out111(conv[111]),.out112(conv[112]),.out113(conv[113]),.out114(conv[114]),.out115(conv[115]),.out116(conv[116]),.out117(conv[117]),.out118(conv[118]),.out119(conv[119]),.out120(conv[120]),.out121(conv[121]),.out122(conv[122]),.out123(conv[123]),.out124(conv[124]),.out125(conv[125]),.out126(conv[126]),.out127(conv[127]),.out128(conv[128]),.out129(conv[129]),.out130(conv[130]),.out131(conv[131]),.out132(conv[132]),.out133(conv[133]),.out134(conv[134]),.out135(conv[135]),.out136(conv[136]),.out137(conv[137]),.out138(conv[138]),.out139(conv[139]),.out140(conv[140]),.out141(conv[141]),.out142(conv[142]),.out143(conv[143]),
.in0(in[0]),.in1(in[1]),.in2(in[2]),.in3(in[3]),.in4(in[4]),.in5(in[5]),.in6(in[6]),.in7(in[7]),.in8(in[8]),.in9(in[9]),.in10(in[10]),.in11(in[11]),.in12(in[12]),.in13(in[13]),.in14(in[14]),.in15(in[15]),.in16(in[16]),.in17(in[17]),.in18(in[18]),.in19(in[19]),.in20(in[20]),.in21(in[21]),.in22(in[22]),.in23(in[23]),.in24(in[24]),.in25(in[25]),.in26(in[26]),.in27(in[27]),.in28(in[28]),.in29(in[29]),.in30(in[30]),.in31(in[31]),.in32(in[32]),.in33(in[33]),.in34(in[34]),.in35(in[35]),.in36(in[36]),.in37(in[37]),.in38(in[38]),.in39(in[39]),.in40(in[40]),.in41(in[41]),.in42(in[42]),.in43(in[43]),.in44(in[44]),.in45(in[45]),.in46(in[46]),.in47(in[47]),.in48(in[48]),.in49(in[49]),.in50(in[50]),.in51(in[51]),.in52(in[52]),.in53(in[53]),.in54(in[54]),.in55(in[55]),.in56(in[56]),.in57(in[57]),.in58(in[58]),.in59(in[59]),.in60(in[60]),.in61(in[61]),.in62(in[62]),.in63(in[63]),.in64(in[64]),.in65(in[65]),.in66(in[66]),.in67(in[67]),.in68(in[68]),.in69(in[69]),.in70(in[70]),.in71(in[71]),.in72(in[72]),.in73(in[73]),.in74(in[74]),.in75(in[75]),.in76(in[76]),.in77(in[77]),.in78(in[78]),.in79(in[79]),.in80(in[80]),.in81(in[81]),.in82(in[82]),.in83(in[83]),.in84(in[84]),.in85(in[85]),.in86(in[86]),.in87(in[87]),.in88(in[88]),.in89(in[89]),.in90(in[90]),.in91(in[91]),.in92(in[92]),.in93(in[93]),.in94(in[94]),.in95(in[95]),.in96(in[96]),.in97(in[97]),.in98(in[98]),.in99(in[99]),.in100(in[100]),.in101(in[101]),.in102(in[102]),.in103(in[103]),.in104(in[104]),.in105(in[105]),.in106(in[106]),.in107(in[107]),.in108(in[108]),.in109(in[109]),.in110(in[110]),.in111(in[111]),.in112(in[112]),.in113(in[113]),.in114(in[114]),.in115(in[115]),.in116(in[116]),.in117(in[117]),.in118(in[118]),.in119(in[119]),.in120(in[120]),.in121(in[121]),.in122(in[122]),.in123(in[123]),.in124(in[124]),.in125(in[125]),.in126(in[126]),.in127(in[127]),.in128(in[128]),.in129(in[129]),.in130(in[130]),.in131(in[131]),.in132(in[132]),.in133(in[133]),.in134(in[134]),.in135(in[135]),.in136(in[136]),.in137(in[137]),.in138(in[138]),.in139(in[139]),.in140(in[140]),.in141(in[141]),.in142(in[142]),.in143(in[143]),.in144(in[144]),.in145(in[145]),.in146(in[146]),.in147(in[147]),.in148(in[148]),.in149(in[149]),.in150(in[150]),.in151(in[151]),.in152(in[152]),.in153(in[153]),.in154(in[154]),.in155(in[155]),.in156(in[156]),.in157(in[157]),.in158(in[158]),.in159(in[159]),.in160(in[160]),.in161(in[161]),.in162(in[162]),.in163(in[163]),.in164(in[164]),.in165(in[165]),.in166(in[166]),.in167(in[167]),.in168(in[168]),.in169(in[169]),.in170(in[170]),.in171(in[171]),.in172(in[172]),.in173(in[173]),.in174(in[174]),.in175(in[175]),.in176(in[176]),.in177(in[177]),.in178(in[178]),.in179(in[179]),.in180(in[180]),.in181(in[181]),.in182(in[182]),.in183(in[183]),.in184(in[184]),.in185(in[185]),.in186(in[186]),.in187(in[187]),.in188(in[188]),.in189(in[189]),.in190(in[190]),.in191(in[191]),.in192(in[192]),.in193(in[193]),.in194(in[194]),.in195(in[195]),.in196(in[196]),.in197(in[197]),.in198(in[198]),.in199(in[199]),.in200(in[200]),.in201(in[201]),.in202(in[202]),.in203(in[203]),.in204(in[204]),.in205(in[205]),.in206(in[206]),.in207(in[207]),.in208(in[208]),.in209(in[209]),.in210(in[210]),.in211(in[211]),.in212(in[212]),.in213(in[213]),.in214(in[214]),.in215(in[215]),.in216(in[216]),.in217(in[217]),.in218(in[218]),.in219(in[219]),.in220(in[220]),.in221(in[221]),.in222(in[222]),.in223(in[223]),.in224(in[224]),.in225(in[225]),.in226(in[226]),.in227(in[227]),.in228(in[228]),.in229(in[229]),.in230(in[230]),.in231(in[231]),.in232(in[232]),.in233(in[233]),.in234(in[234]),.in235(in[235]),.in236(in[236]),.in237(in[237]),.in238(in[238]),.in239(in[239]),.in240(in[240]),.in241(in[241]),.in242(in[242]),.in243(in[243]),.in244(in[244]),.in245(in[245]),.in246(in[246]),.in247(in[247]),.in248(in[248]),.in249(in[249]),.in250(in[250]),.in251(in[251]),.in252(in[252]),.in253(in[253]),.in254(in[254]),.in255(in[255]),.in256(in[256]),.in257(in[257]),.in258(in[258]),.in259(in[259]),.in260(in[260]),.in261(in[261]),.in262(in[262]),.in263(in[263]),.in264(in[264]),.in265(in[265]),.in266(in[266]),.in267(in[267]),.in268(in[268]),.in269(in[269]),.in270(in[270]),.in271(in[271]),.in272(in[272]),.in273(in[273]),.in274(in[274]),.in275(in[275]),.in276(in[276]),.in277(in[277]),.in278(in[278]),.in279(in[279]),.in280(in[280]),.in281(in[281]),.in282(in[282]),.in283(in[283]),.in284(in[284]),.in285(in[285]),.in286(in[286]),.in287(in[287]),.in288(in[288]),.in289(in[289]),.in290(in[290]),.in291(in[291]),.in292(in[292]),.in293(in[293]),.in294(in[294]),.in295(in[295]),.in296(in[296]),.in297(in[297]),.in298(in[298]),.in299(in[299]),.in300(in[300]),.in301(in[301]),.in302(in[302]),.in303(in[303]),.in304(in[304]),.in305(in[305]),.in306(in[306]),.in307(in[307]),.in308(in[308]),.in309(in[309]),.in310(in[310]),.in311(in[311]),.in312(in[312]),.in313(in[313]),.in314(in[314]),.in315(in[315]),.in316(in[316]),.in317(in[317]),.in318(in[318]),.in319(in[319]),.in320(in[320]),.in321(in[321]),.in322(in[322]),.in323(in[323]),.in324(in[324]),.in325(in[325]),.in326(in[326]),.in327(in[327]),.in328(in[328]),.in329(in[329]),.in330(in[330]),.in331(in[331]),.in332(in[332]),.in333(in[333]),.in334(in[334]),.in335(in[335]),.in336(in[336]),.in337(in[337]),.in338(in[338]),.in339(in[339]),.in340(in[340]),.in341(in[341]),.in342(in[342]),.in343(in[343]),.in344(in[344]),.in345(in[345]),.in346(in[346]),.in347(in[347]),.in348(in[348]),.in349(in[349]),.in350(in[350]),.in351(in[351]),.in352(in[352]),.in353(in[353]),.in354(in[354]),.in355(in[355]),.in356(in[356]),.in357(in[357]),.in358(in[358]),.in359(in[359]),.in360(in[360]),.in361(in[361]),.in362(in[362]),.in363(in[363]),.in364(in[364]),.in365(in[365]),.in366(in[366]),.in367(in[367]),.in368(in[368]),.in369(in[369]),.in370(in[370]),.in371(in[371]),.in372(in[372]),.in373(in[373]),.in374(in[374]),.in375(in[375]),.in376(in[376]),.in377(in[377]),.in378(in[378]),.in379(in[379]),.in380(in[380]),.in381(in[381]),.in382(in[382]),.in383(in[383]),.in384(in[384]),.in385(in[385]),.in386(in[386]),.in387(in[387]),.in388(in[388]),.in389(in[389]),.in390(in[390]),.in391(in[391]),.in392(in[392]),.in393(in[393]),.in394(in[394]),.in395(in[395]),.in396(in[396]),.in397(in[397]),.in398(in[398]),.in399(in[399]),.in400(in[400]),.in401(in[401]),.in402(in[402]),.in403(in[403]),.in404(in[404]),.in405(in[405]),.in406(in[406]),.in407(in[407]),.in408(in[408]),.in409(in[409]),.in410(in[410]),.in411(in[411]),.in412(in[412]),.in413(in[413]),.in414(in[414]),.in415(in[415]),.in416(in[416]),.in417(in[417]),.in418(in[418]),.in419(in[419]),.in420(in[420]),.in421(in[421]),.in422(in[422]),.in423(in[423]),.in424(in[424]),.in425(in[425]),.in426(in[426]),.in427(in[427]),.in428(in[428]),.in429(in[429]),.in430(in[430]),.in431(in[431]),.in432(in[432]),.in433(in[433]),.in434(in[434]),.in435(in[435]),.in436(in[436]),.in437(in[437]),.in438(in[438]),.in439(in[439]),.in440(in[440]),.in441(in[441]),.in442(in[442]),.in443(in[443]),.in444(in[444]),.in445(in[445]),.in446(in[446]),.in447(in[447]),.in448(in[448]),.in449(in[449]),.in450(in[450]),.in451(in[451]),.in452(in[452]),.in453(in[453]),.in454(in[454]),.in455(in[455]),.in456(in[456]),.in457(in[457]),.in458(in[458]),.in459(in[459]),.in460(in[460]),.in461(in[461]),.in462(in[462]),.in463(in[463]),.in464(in[464]),.in465(in[465]),.in466(in[466]),.in467(in[467]),.in468(in[468]),.in469(in[469]),.in470(in[470]),.in471(in[471]),.in472(in[472]),.in473(in[473]),.in474(in[474]),.in475(in[475]),.in476(in[476]),.in477(in[477]),.in478(in[478]),.in479(in[479]),.in480(in[480]),.in481(in[481]),.in482(in[482]),.in483(in[483]),.in484(in[484]),.in485(in[485]),.in486(in[486]),.in487(in[487]),.in488(in[488]),.in489(in[489]),.in490(in[490]),.in491(in[491]),.in492(in[492]),.in493(in[493]),.in494(in[494]),.in495(in[495]),.in496(in[496]),.in497(in[497]),.in498(in[498]),.in499(in[499]),.in500(in[500]),.in501(in[501]),.in502(in[502]),.in503(in[503]),.in504(in[504]),.in505(in[505]),.in506(in[506]),.in507(in[507]),.in508(in[508]),.in509(in[509]),.in510(in[510]),.in511(in[511]),.in512(in[512]),.in513(in[513]),.in514(in[514]),.in515(in[515]),.in516(in[516]),.in517(in[517]),.in518(in[518]),.in519(in[519]),.in520(in[520]),.in521(in[521]),.in522(in[522]),.in523(in[523]),.in524(in[524]),.in525(in[525]),.in526(in[526]),.in527(in[527]),.in528(in[528]),.in529(in[529]),.in530(in[530]),.in531(in[531]),.in532(in[532]),.in533(in[533]),.in534(in[534]),.in535(in[535]),.in536(in[536]),.in537(in[537]),.in538(in[538]),.in539(in[539]),.in540(in[540]),.in541(in[541]),.in542(in[542]),.in543(in[543]),.in544(in[544]),.in545(in[545]),.in546(in[546]),.in547(in[547]),.in548(in[548]),.in549(in[549]),.in550(in[550]),.in551(in[551]),.in552(in[552]),.in553(in[553]),.in554(in[554]),.in555(in[555]),.in556(in[556]),.in557(in[557]),.in558(in[558]),.in559(in[559]),.in560(in[560]),.in561(in[561]),.in562(in[562]),.in563(in[563]),.in564(in[564]),.in565(in[565]),.in566(in[566]),.in567(in[567]),.in568(in[568]),.in569(in[569]),.in570(in[570]),.in571(in[571]),.in572(in[572]),.in573(in[573]),.in574(in[574]),.in575(in[575]),
.clk(clk),.ready(ready),.start(start));*/

/*ConvLayer ConvLayer1(.ready(ready),.weight0(weight[0]), .weight1(weight[1]), .weight2(weight[2]), .weight3(weight[3]),.weight4(weight[4]), .weight5(weight[5]), .weight6(weight[6]), .weight7(weight[7]),.weight8(weight[8]), .weight9(weight[9]), .weight10(weight[10]), .weight11(weight[11]), .weight12(weight[12]),.weight13(weight[13]), .weight14(weight[14]), .weight15(weight[15]), .weight16(weight[16]), .weight17(weight[17]), .weight18(weight[18]), .weight19(weight[19]), .weight20(weight[20]), .weight21(weight[21]), .weight22(weight[22]), .weight23(weight[23]), .weight24(weight[24]),.in0(in[0]),.in1(in[1]),.in2(in[2]),.in3(in[3]),.in4(in[4]),.in5(in[5]),.in6(in[6]),.in7(in[7]),.in8(in[8]),.in9(in[9]),.in10(in[10]),.in11(in[11]),.in12(in[12]),.in13(in[13]),.in14(in[14]),.in15(in[15]),.in16(in[16]),.in17(in[17]),.in18(in[18]),.in19(in[19]),.in20(in[20]),.in21(in[21]),.in22(in[22]),.in23(in[23]),.in24(in[24]),.in25(in[25]),.in26(in[26]),.in27(in[27]),.in28(in[28]),.in29(in[29]),.in30(in[30]),.in31(in[31]),.in32(in[32]),.in33(in[33]),.in34(in[34]),.in35(in[35]),.in36(in[36]),.in37(in[37]),.in38(in[38]),.in39(in[39]),.in40(in[40]),.in41(in[41]),.in42(in[42]),.in43(in[43]),.in44(in[44]),.in45(in[45]),.in46(in[46]),.in47(in[47]),.in48(in[48]),.in49(in[49]),.in50(in[50]),.in51(in[51]),.in52(in[52]),.in53(in[53]),.in54(in[54]),.in55(in[55]),.in56(in[56]),.in57(in[57]),.in58(in[58]),.in59(in[59]),.in60(in[60]),.in61(in[61]),.in62(in[62]),.in63(in[63]),.in64(in[64]),.in65(in[65]),.in66(in[66]),.in67(in[67]),.in68(in[68]),.in69(in[69]),.in70(in[70]),.in71(in[71]),.in72(in[72]),.in73(in[73]),.in74(in[74]),.in75(in[75]),.in76(in[76]),.in77(in[77]),.in78(in[78]),.in79(in[79]),
.in80(in[80]),.in81(in[81]),.in82(in[82]),.in83(in[83]),.in84(in[84]),.in85(in[85]),.in86(in[86]),.in87(in[87]),.in88(in[88]),.in89(in[89]),.in90(in[90]),.in91(in[91]),.in92(in[92]),.in93(in[93]),.in94(in[94]),.in95(in[95]),.in96(in[96]),.in97(in[97]),.in98(in[98]),.in99(in[99]),.in100(in[100]),.in101(in[101]),.in102(in[102]),.in103(in[103]),.in104(in[104]),.in105(in[105]),.in106(in[106]),.in107(in[107]),.in108(in[108]),.in109(in[109]),.in110(in[110]),.in111(in[111]),.in112(in[112]),.in113(in[113]),.in114(in[114]),.in115(in[115]),.in116(in[116]),.in117(in[117]),.in118(in[118]),.in119(in[119]),.in120(in[120]),.in121(in[121]),.in122(in[122]),.in123(in[123]),.in124(in[124]),.in125(in[125]),.in126(in[126]),.in127(in[127]),.in128(in[128]),.in129(in[129]),.in130(in[130]),.in131(in[131]),.in132(in[132]),.in133(in[133]),.in134(in[134]),.in135(in[135]),.in136(in[136]),.in137(in[137]),.in138(in[138]),.in139(in[139]),.in140(in[140]),.in141(in[141]),.in142(in[142]),.in143(in[143]),.in144(in[144]),.in145(in[145]),.in146(in[146]),.in147(in[147]),.in148(in[148]),.in149(in[149]),.in150(in[150]),.in151(in[151]),.in152(in[152]),.in153(in[153]),.in154(in[154]),.in155(in[155]),.in156(in[156]),.in157(in[157]),.in158(in[158]),.in159(in[159]),.in160(in[160]),.in161(in[161]),.in162(in[162]),.in163(in[163]),.in164(in[164]),.in165(in[165]),.in166(in[166]),.in167(in[167]),.in168(in[168]),.in169(in[169]),.in170(in[170]),.in171(in[171]),.in172(in[172]),.in173(in[173]),.in174(in[174]),.in175(in[175]),.in176(in[176]),.in177(in[177]),.in178(in[178]),.in179(in[179]),.in180(in[180]),.in181(in[181]),.in182(in[182]),.in183(in[183]),.in184(in[184]),.in185(in[185]),.in186(in[186]),.in187(in[187]),.in188(in[188]),.in189(in[189]),.in190(in[190]),.in191(in[191]),.in192(in[192]),.in193(in[193]),.in194(in[194]),.in195(in[195]),.in196(in[196]),.in197(in[197]),.in198(in[198]),.in199(in[199]),.in200(in[200]),.in201(in[201]),.in202(in[202]),.in203(in[203]),.in204(in[204]),.in205(in[205]),.in206(in[206]),.in207(in[207]),.in208(in[208]),.in209(in[209]),.in210(in[210]),.in211(in[211]),.in212(in[212]),.in213(in[213]),.in214(in[214]),.in215(in[215]),.in216(in[216]),.in217(in[217]),.in218(in[218]),.in219(in[219]),.in220(in[220]),.in221(in[221]),.in222(in[222]),.in223(in[223]),.in224(in[224]),.in225(in[225]),.in226(in[226]),.in227(in[227]),.in228(in[228]),.in229(in[229]),.in230(in[230]),.in231(in[231]),.in232(in[232]),.in233(in[233]),.in234(in[234]),.in235(in[235]),.in236(in[236]),.in237(in[237]),.in238(in[238]),.in239(in[239]),.in240(in[240]),.in241(in[241]),.in242(in[242]),.in243(in[243]),.in244(in[244]),.in245(in[245]),.in246(in[246]),.in247(in[247]),.in248(in[248]),.in249(in[249]),.in250(in[250]),.in251(in[251]),.in252(in[252]),.in253(in[253]),.in254(in[254]),.in255(in[255]),.in256(in[256]),.in257(in[257]),.in258(in[258]),.in259(in[259]),.in260(in[260]),.in261(in[261]),.in262(in[262]),.in263(in[263]),.in264(in[264]),.in265(in[265]),.in266(in[266]),.in267(in[267]),.in268(in[268]),.in269(in[269]),.in270(in[270]),.in271(in[271]),.in272(in[272]),.in273(in[273]),.in274(in[274]),.in275(in[275]),.in276(in[276]),.in277(in[277]),.in278(in[278]),.in279(in[279]),.in280(in[280]),.in281(in[281]),.in282(in[282]),.in283(in[283]),.in284(in[284]),.in285(in[285]),.in286(in[286]),.in287(in[287]),.in288(in[288]),.in289(in[289]),.in290(in[290]),.in291(in[291]),.in292(in[292]),.in293(in[293]),.in294(in[294]),.in295(in[295]),.in296(in[296]),.in297(in[297]),.in298(in[298]),.in299(in[299]),.in300(in[300]),.in301(in[301]),.in302(in[302]),.in303(in[303]),.in304(in[304]),.in305(in[305]),.in306(in[306]),.in307(in[307]),.in308(in[308]),.in309(in[309]),.in310(in[310]),.in311(in[311]),.in312(in[312]),.in313(in[313]),.in314(in[314]),.in315(in[315]),.in316(in[316]),.in317(in[317]),.in318(in[318]),.in319(in[319]),.in320(in[320]),.in321(in[321]),.in322(in[322]),.in323(in[323]),.in324(in[324]),.in325(in[325]),.in326(in[326]),.in327(in[327]),.in328(in[328]),.in329(in[329]),.in330(in[330]),.in331(in[331]),.in332(in[332]),.in333(in[333]),.in334(in[334]),.in335(in[335]),.in336(in[336]),.in337(in[337]),.in338(in[338]),.in339(in[339]),.in340(in[340]),.in341(in[341]),.in342(in[342]),.in343(in[343]),.in344(in[344]),.in345(in[345]),.in346(in[346]),.in347(in[347]),.in348(in[348]),.in349(in[349]),.in350(in[350]),.in351(in[351]),.in352(in[352]),.in353(in[353]),.in354(in[354]),.in355(in[355]),.in356(in[356]),.in357(in[357]),.in358(in[358]),.in359(in[359]),.in360(in[360]),.in361(in[361]),.in362(in[362]),.in363(in[363]),.in364(in[364]),.in365(in[365]),.in366(in[366]),.in367(in[367]),.in368(in[368]),.in369(in[369]),.in370(in[370]),.in371(in[371]),.in372(in[372]),.in373(in[373]),.in374(in[374]),.in375(in[375]),.in376(in[376]),.in377(in[377]),.in378(in[378]),.in379(in[379]),.in380(in[380]),.in381(in[381]),.in382(in[382]),.in383(in[383]),.in384(in[384]),.in385(in[385]),.in386(in[386]),.in387(in[387]),.in388(in[388]),.in389(in[389]),.in390(in[390]),.in391(in[391]),.in392(in[392]),.in393(in[393]),.in394(in[394]),.in395(in[395]),.in396(in[396]),.in397(in[397]),.in398(in[398]),.in399(in[399]),.in400(in[400]),.in401(in[401]),.in402(in[402]),.in403(in[403]),.in404(in[404]),.in405(in[405]),.in406(in[406]),.in407(in[407]),.in408(in[408]),.in409(in[409]),.in410(in[410]),.in411(in[411]),.in412(in[412]),.in413(in[413]),.in414(in[414]),.in415(in[415]),.in416(in[416]),.in417(in[417]),.in418(in[418]),.in419(in[419]),.in420(in[420]),.in421(in[421]),.in422(in[422]),.in423(in[423]),.in424(in[424]),.in425(in[425]),.in426(in[426]),.in427(in[427]),.in428(in[428]),.in429(in[429]),.in430(in[430]),.in431(in[431]),.in432(in[432]),.in433(in[433]),.in434(in[434]),.in435(in[435]),.in436(in[436]),.in437(in[437]),.in438(in[438]),.in439(in[439]),.in440(in[440]),.in441(in[441]),.in442(in[442]),.in443(in[443]),.in444(in[444]),.in445(in[445]),.in446(in[446]),.in447(in[447]),.in448(in[448]),.in449(in[449]),.in450(in[450]),.in451(in[451]),.in452(in[452]),.in453(in[453]),.in454(in[454]),.in455(in[455]),.in456(in[456]),.in457(in[457]),.in458(in[458]),.in459(in[459]),.in460(in[460]),.in461(in[461]),.in462(in[462]),.in463(in[463]),.in464(in[464]),.in465(in[465]),.in466(in[466]),.in467(in[467]),.in468(in[468]),.in469(in[469]),.in470(in[470]),.in471(in[471]),.in472(in[472]),.in473(in[473]),.in474(in[474]),.in475(in[475]),.in476(in[476]),.in477(in[477]),.in478(in[478]),.in479(in[479]),.in480(in[480]),.in481(in[481]),.in482(in[482]),.in483(in[483]),.in484(in[484]),.in485(in[485]),.in486(in[486]),.in487(in[487]),.in488(in[488]),.in489(in[489]),.in490(in[490]),.in491(in[491]),.in492(in[492]),.in493(in[493]),.in494(in[494]),.in495(in[495]),.in496(in[496]),.in497(in[497]),.in498(in[498]),.in499(in[499]),.in500(in[500]),.in501(in[501]),.in502(in[502]),.in503(in[503]),.in504(in[504]),.in505(in[505]),.in506(in[506]),.in507(in[507]),.in508(in[508]),.in509(in[509]),.in510(in[510]),.in511(in[511]),.in512(in[512]),.in513(in[513]),.in514(in[514]),.in515(in[515]),.in516(in[516]),.in517(in[517]),.in518(in[518]),.in519(in[519]),.in520(in[520]),.in521(in[521]),.in522(in[522]),.in523(in[523]),.in524(in[524]),.in525(in[525]),.in526(in[526]),.in527(in[527]),.in528(in[528]),.in529(in[529]),.in530(in[530]),.in531(in[531]),.in532(in[532]),.in533(in[533]),.in534(in[534]),.in535(in[535]),.in536(in[536]),.in537(in[537]),.in538(in[538]),.in539(in[539]),.in540(in[540]),.in541(in[541]),.in542(in[542]),.in543(in[543]),.in544(in[544]),.in545(in[545]),.in546(in[546]),.in547(in[547]),.in548(in[548]),.in549(in[549]),.in550(in[550]),.in551(in[551]),.in552(in[552]),.in553(in[553]),.in554(in[554]),.in555(in[555]),.in556(in[556]),.in557(in[557]),.in558(in[558]),.in559(in[559]),.in560(in[560]),.in561(in[561]),.in562(in[562]),.in563(in[563]),.in564(in[564]),.in565(in[565]),.in566(in[566]),.in567(in[567]),.in568(in[568]),.in569(in[569]),.in570(in[570]),.in571(in[571]),.in572(in[572]),.in573(in[573]),.in574(in[574]),.in575(in[575]),.in576(in[576]),.in577(in[577]),.in578(in[578]),.in579(in[579]),.in580(in[580]),.in581(in[581]),.in582(in[582]),.in583(in[583]),.in584(in[584]),.in585(in[585]),.in586(in[586]),.in587(in[587]),.in588(in[588]),.in589(in[589]),.in590(in[590]),.in591(in[591]),.in592(in[592]),.in593(in[593]),.in594(in[594]),.in595(in[595]),.in596(in[596]),.in597(in[597]),.in598(in[598]),.in599(in[599]),.in600(in[600]),.in601(in[601]),.in602(in[602]),.in603(in[603]),.in604(in[604]),.in605(in[605]),.in606(in[606]),.in607(in[607]),.in608(in[608]),.in609(in[609]),.in610(in[610]),.in611(in[611]),.in612(in[612]),.in613(in[613]),.in614(in[614]),.in615(in[615]),.in616(in[616]),.in617(in[617]),.in618(in[618]),.in619(in[619]),.in620(in[620]),.in621(in[621]),.in622(in[622]),.in623(in[623]),.in624(in[624]),.in625(in[625]),.in626(in[626]),.in627(in[627]),.in628(in[628]),.in629(in[629]),.in630(in[630]),.in631(in[631]),.in632(in[632]),.in633(in[633]),.in634(in[634]),.in635(in[635]),.in636(in[636]),.in637(in[637]),.in638(in[638]),.in639(in[639]),.in640(in[640]),.in641(in[641]),.in642(in[642]),.in643(in[643]),.in644(in[644]),.in645(in[645]),.in646(in[646]),.in647(in[647]),.in648(in[648]),.in649(in[649]),.in650(in[650]),.in651(in[651]),.in652(in[652]),.in653(in[653]),.in654(in[654]),.in655(in[655]),.in656(in[656]),.in657(in[657]),.in658(in[658]),.in659(in[659]),.in660(in[660]),.in661(in[661]),.in662(in[662]),.in663(in[663]),.in664(in[664]),.in665(in[665]),.in666(in[666]),.in667(in[667]),.in668(in[668]),.in669(in[669]),.in670(in[670]),.in671(in[671]),.in672(in[672]),.in673(in[673]),.in674(in[674]),.in675(in[675]),.in676(in[676]),.in677(in[677]),.in678(in[678]),.in679(in[679]),.in680(in[680]),.in681(in[681]),.in682(in[682]),.in683(in[683]),.in684(in[684]),.in685(in[685]),.in686(in[686]),.in687(in[687]),.in688(in[688]),.in689(in[689]),.in690(in[690]),.in691(in[691]),.in692(in[692]),.in693(in[693]),.in694(in[694]),.in695(in[695]),.in696(in[696]),.in697(in[697]),.in698(in[698]),.in699(in[699]),.in700(in[700]),.in701(in[701]),.in702(in[702]),.in703(in[703]),.in704(in[704]),.in705(in[705]),.in706(in[706]),.in707(in[707]),.in708(in[708]),.in709(in[709]),.in710(in[710]),.in711(in[711]),.in712(in[712]),.in713(in[713]),.in714(in[714]),.in715(in[715]),.in716(in[716]),.in717(in[717]),.in718(in[718]),.in719(in[719]),.in720(in[720]),.in721(in[721]),.in722(in[722]),.in723(in[723]),.in724(in[724]),.in725(in[725]),.in726(in[726]),.in727(in[727]),.in728(in[728]),.in729(in[729]),.in730(in[730]),.in731(in[731]),.in732(in[732]),.in733(in[733]),.in734(in[734]),.in735(in[735]),.in736(in[736]),.in737(in[737]),.in738(in[738]),.in739(in[739]),.in740(in[740]),.in741(in[741]),.in742(in[742]),.in743(in[743]),.in744(in[744]),.in745(in[745]),.in746(in[746]),.in747(in[747]),.in748(in[748]),.in749(in[749]),.in750(in[750]),.in751(in[751]),.in752(in[752]),.in753(in[753]),.in754(in[754]),.in755(in[755]),.in756(in[756]),.in757(in[757]),.in758(in[758]),.in759(in[759]),.in760(in[760]),.in761(in[761]),.in762(in[762]),.in763(in[763]),.in764(in[764]),.in765(in[765]),.in766(in[766]),.in767(in[767]),.in768(in[768]),.in769(in[769]),.in770(in[770]),.in771(in[771]),.in772(in[772]),.in773(in[773]),.in774(in[774]),.in775(in[775]),.in776(in[776]),.in777(in[777]),.in778(in[778]),.in779(in[779]),.in780(in[780]),.in781(in[781]),.in782(in[782]),.in783(in[783]),.bias(bias), .clk(clk),.conv0(conv[0]),.conv1(conv[1]),.conv2(conv[2]),.conv3(conv[3]),.conv4(conv[4]),.conv5(conv[5]),.conv6(conv[6]),.conv7(conv[7]),.conv8(conv[8]),.conv9(conv[9]),.conv10(conv[10]),.conv11(conv[11]),.conv12(conv[12]),.conv13(conv[13]),.conv14(conv[14]),.conv15(conv[15]),.conv16(conv[16]),.conv17(conv[17]),.conv18(conv[18]),.conv19(conv[19]),.conv20(conv[20]),.conv21(conv[21]),.conv22(conv[22]),.conv23(conv[23]),.conv24(conv[24]),.conv25(conv[25]),.conv26(conv[26]),.conv27(conv[27]),.conv28(conv[28]),.conv29(conv[29]),.conv30(conv[30]),.conv31(conv[31]),.conv32(conv[32]),.conv33(conv[33]),.conv34(conv[34]),.conv35(conv[35]),.conv36(conv[36]),.conv37(conv[37]),.conv38(conv[38]),.conv39(conv[39]),.conv40(conv[40]),.conv41(conv[41]),.conv42(conv[42]),.conv43(conv[43]),.conv44(conv[44]),.conv45(conv[45]),.conv46(conv[46]),.conv47(conv[47]),.conv48(conv[48]),.conv49(conv[49]),.conv50(conv[50]),.conv51(conv[51]),.conv52(conv[52]),.conv53(conv[53]),.conv54(conv[54]),.conv55(conv[55]),.conv56(conv[56]),.conv57(conv[57]),.conv58(conv[58]),.conv59(conv[59]),.conv60(conv[60]),.conv61(conv[61]),.conv62(conv[62]),.conv63(conv[63]),.conv64(conv[64]),.conv65(conv[65]),.conv66(conv[66]),.conv67(conv[67]),.conv68(conv[68]),.conv69(conv[69]),.conv70(conv[70]),.conv71(conv[71]),.conv72(conv[72]),.conv73(conv[73]),.conv74(conv[74]),.conv75(conv[75]),.conv76(conv[76]),.conv77(conv[77]),.conv78(conv[78]),.conv79(conv[79]),.conv80(conv[80]),.conv81(conv[81]),.conv82(conv[82]),.conv83(conv[83]),.conv84(conv[84]),.conv85(conv[85]),.conv86(conv[86]),.conv87(conv[87]),.conv88(conv[88]),.conv89(conv[89]),.conv90(conv[90]),.conv91(conv[91]),.conv92(conv[92]),.conv93(conv[93]),.conv94(conv[94]),.conv95(conv[95]),.conv96(conv[96]),.conv97(conv[97]),.conv98(conv[98]),.conv99(conv[99]),.conv100(conv[100]),.conv101(conv[101]),.conv102(conv[102]),.conv103(conv[103]),.conv104(conv[104]),.conv105(conv[105]),.conv106(conv[106]),.conv107(conv[107]),.conv108(conv[108]),.conv109(conv[109]),.conv110(conv[110]),.conv111(conv[111]),.conv112(conv[112]),.conv113(conv[113]),.conv114(conv[114]),.conv115(conv[115]),.conv116(conv[116]),.conv117(conv[117]),.conv118(conv[118]),.conv119(conv[119]),.conv120(conv[120]),.conv121(conv[121]),.conv122(conv[122]),.conv123(conv[123]),.conv124(conv[124]),.conv125(conv[125]),.conv126(conv[126]),.conv127(conv[127]),.conv128(conv[128]),.conv129(conv[129]),.conv130(conv[130]),.conv131(conv[131]),.conv132(conv[132]),.conv133(conv[133]),.conv134(conv[134]),.conv135(conv[135]),.conv136(conv[136]),.conv137(conv[137]),.conv138(conv[138]),.conv139(conv[139]),.conv140(conv[140]),.conv141(conv[141]),.conv142(conv[142]),.conv143(conv[143]),.conv144(conv[144]),.conv145(conv[145]),.conv146(conv[146]),.conv147(conv[147]),.conv148(conv[148]),.conv149(conv[149]),.conv150(conv[150]),.conv151(conv[151]),.conv152(conv[152]),.conv153(conv[153]),.conv154(conv[154]),.conv155(conv[155]),.conv156(conv[156]),.conv157(conv[157]),.conv158(conv[158]),.conv159(conv[159]),.conv160(conv[160]),.conv161(conv[161]),.conv162(conv[162]),.conv163(conv[163]),.conv164(conv[164]),.conv165(conv[165]),.conv166(conv[166]),.conv167(conv[167]),.conv168(conv[168]),.conv169(conv[169]),.conv170(conv[170]),.conv171(conv[171]),.conv172(conv[172]),.conv173(conv[173]),.conv174(conv[174]),.conv175(conv[175]),.conv176(conv[176]),.conv177(conv[177]),.conv178(conv[178]),.conv179(conv[179]),.conv180(conv[180]),.conv181(conv[181]),.conv182(conv[182]),.conv183(conv[183]),.conv184(conv[184]),.conv185(conv[185]),.conv186(conv[186]),.conv187(conv[187]),.conv188(conv[188]),.conv189(conv[189]),.conv190(conv[190]),.conv191(conv[191]),.conv192(conv[192]),.conv193(conv[193]),.conv194(conv[194]),.conv195(conv[195]),.conv196(conv[196]),.conv197(conv[197]),.conv198(conv[198]),.conv199(conv[199]),.conv200(conv[200]),.conv201(conv[201]),.conv202(conv[202]),.conv203(conv[203]),.conv204(conv[204]),.conv205(conv[205]),.conv206(conv[206]),.conv207(conv[207]),.conv208(conv[208]),.conv209(conv[209]),.conv210(conv[210]),.conv211(conv[211]),.conv212(conv[212]),.conv213(conv[213]),.conv214(conv[214]),.conv215(conv[215]),.conv216(conv[216]),.conv217(conv[217]),.conv218(conv[218]),.conv219(conv[219]),.conv220(conv[220]),.conv221(conv[221]),.conv222(conv[222]),.conv223(conv[223]),.conv224(conv[224]),.conv225(conv[225]),.conv226(conv[226]),.conv227(conv[227]),.conv228(conv[228]),.conv229(conv[229]),.conv230(conv[230]),.conv231(conv[231]),.conv232(conv[232]),.conv233(conv[233]),.conv234(conv[234]),.conv235(conv[235]),.conv236(conv[236]),.conv237(conv[237]),.conv238(conv[238]),.conv239(conv[239]),.conv240(conv[240]),.conv241(conv[241]),.conv242(conv[242]),.conv243(conv[243]),.conv244(conv[244]),.conv245(conv[245]),.conv246(conv[246]),.conv247(conv[247]),.conv248(conv[248]),.conv249(conv[249]),.conv250(conv[250]),.conv251(conv[251]),.conv252(conv[252]),.conv253(conv[253]),.conv254(conv[254]),.conv255(conv[255]),.conv256(conv[256]),.conv257(conv[257]),.conv258(conv[258]),.conv259(conv[259]),.conv260(conv[260]),.conv261(conv[261]),.conv262(conv[262]),.conv263(conv[263]),.conv264(conv[264]),.conv265(conv[265]),.conv266(conv[266]),.conv267(conv[267]),.conv268(conv[268]),.conv269(conv[269]),.conv270(conv[270]),.conv271(conv[271]),.conv272(conv[272]),.conv273(conv[273]),.conv274(conv[274]),.conv275(conv[275]),.conv276(conv[276]),.conv277(conv[277]),.conv278(conv[278]),.conv279(conv[279]),.conv280(conv[280]),.conv281(conv[281]),.conv282(conv[282]),.conv283(conv[283]),.conv284(conv[284]),.conv285(conv[285]),.conv286(conv[286]),.conv287(conv[287]),.conv288(conv[288]),.conv289(conv[289]),.conv290(conv[290]),.conv291(conv[291]),.conv292(conv[292]),.conv293(conv[293]),.conv294(conv[294]),.conv295(conv[295]),.conv296(conv[296]),.conv297(conv[297]),.conv298(conv[298]),.conv299(conv[299]),.conv300(conv[300]),.conv301(conv[301]),.conv302(conv[302]),.conv303(conv[303]),.conv304(conv[304]),.conv305(conv[305]),.conv306(conv[306]),.conv307(conv[307]),.conv308(conv[308]),.conv309(conv[309]),.conv310(conv[310]),.conv311(conv[311]),.conv312(conv[312]),.conv313(conv[313]),.conv314(conv[314]),.conv315(conv[315]),.conv316(conv[316]),.conv317(conv[317]),.conv318(conv[318]),.conv319(conv[319]),.conv320(conv[320]),.conv321(conv[321]),.conv322(conv[322]),.conv323(conv[323]),.conv324(conv[324]),.conv325(conv[325]),.conv326(conv[326]),.conv327(conv[327]),.conv328(conv[328]),.conv329(conv[329]),.conv330(conv[330]),.conv331(conv[331]),.conv332(conv[332]),.conv333(conv[333]),.conv334(conv[334]),.conv335(conv[335]),.conv336(conv[336]),.conv337(conv[337]),.conv338(conv[338]),.conv339(conv[339]),.conv340(conv[340]),.conv341(conv[341]),.conv342(conv[342]),.conv343(conv[343]),.conv344(conv[344]),.conv345(conv[345]),.conv346(conv[346]),.conv347(conv[347]),.conv348(conv[348]),.conv349(conv[349]),.conv350(conv[350]),.conv351(conv[351]),.conv352(conv[352]),.conv353(conv[353]),.conv354(conv[354]),.conv355(conv[355]),.conv356(conv[356]),.conv357(conv[357]),.conv358(conv[358]),.conv359(conv[359]),.conv360(conv[360]),.conv361(conv[361]),.conv362(conv[362]),.conv363(conv[363]),.conv364(conv[364]),.conv365(conv[365]),.conv366(conv[366]),.conv367(conv[367]),.conv368(conv[368]),.conv369(conv[369]),.conv370(conv[370]),.conv371(conv[371]),.conv372(conv[372]),.conv373(conv[373]),.conv374(conv[374]),.conv375(conv[375]),.conv376(conv[376]),.conv377(conv[377]),.conv378(conv[378]),.conv379(conv[379]),.conv380(conv[380]),.conv381(conv[381]),.conv382(conv[382]),.conv383(conv[383]),.conv384(conv[384]),.conv385(conv[385]),.conv386(conv[386]),.conv387(conv[387]),.conv388(conv[388]),.conv389(conv[389]),.conv390(conv[390]),.conv391(conv[391]),.conv392(conv[392]),.conv393(conv[393]),.conv394(conv[394]),.conv395(conv[395]),.conv396(conv[396]),.conv397(conv[397]),.conv398(conv[398]),.conv399(conv[399]),.conv400(conv[400]),.conv401(conv[401]),.conv402(conv[402]),.conv403(conv[403]),.conv404(conv[404]),.conv405(conv[405]),.conv406(conv[406]),.conv407(conv[407]),.conv408(conv[408]),.conv409(conv[409]),.conv410(conv[410]),.conv411(conv[411]),.conv412(conv[412]),.conv413(conv[413]),.conv414(conv[414]),.conv415(conv[415]),.conv416(conv[416]),.conv417(conv[417]),.conv418(conv[418]),.conv419(conv[419]),.conv420(conv[420]),.conv421(conv[421]),.conv422(conv[422]),.conv423(conv[423]),.conv424(conv[424]),.conv425(conv[425]),.conv426(conv[426]),.conv427(conv[427]),.conv428(conv[428]),.conv429(conv[429]),.conv430(conv[430]),.conv431(conv[431]),.conv432(conv[432]),.conv433(conv[433]),.conv434(conv[434]),.conv435(conv[435]),.conv436(conv[436]),.conv437(conv[437]),.conv438(conv[438]),.conv439(conv[439]),.conv440(conv[440]),.conv441(conv[441]),.conv442(conv[442]),.conv443(conv[443]),.conv444(conv[444]),.conv445(conv[445]),.conv446(conv[446]),.conv447(conv[447]),.conv448(conv[448]),.conv449(conv[449]),.conv450(conv[450]),.conv451(conv[451]),.conv452(conv[452]),.conv453(conv[453]),.conv454(conv[454]),.conv455(conv[455]),.conv456(conv[456]),.conv457(conv[457]),.conv458(conv[458]),.conv459(conv[459]),.conv460(conv[460]),.conv461(conv[461]),.conv462(conv[462]),.conv463(conv[463]),.conv464(conv[464]),.conv465(conv[465]),.conv466(conv[466]),.conv467(conv[467]),.conv468(conv[468]),.conv469(conv[469]),.conv470(conv[470]),.conv471(conv[471]),.conv472(conv[472]),.conv473(conv[473]),.conv474(conv[474]),.conv475(conv[475]),.conv476(conv[476]),.conv477(conv[477]),.conv478(conv[478]),.conv479(conv[479]),.conv480(conv[480]),.conv481(conv[481]),.conv482(conv[482]),.conv483(conv[483]),.conv484(conv[484]),.conv485(conv[485]),.conv486(conv[486]),.conv487(conv[487]),.conv488(conv[488]),.conv489(conv[489]),.conv490(conv[490]),.conv491(conv[491]),.conv492(conv[492]),.conv493(conv[493]),.conv494(conv[494]),.conv495(conv[495]),.conv496(conv[496]),.conv497(conv[497]),.conv498(conv[498]),.conv499(conv[499]),.conv500(conv[500]),.conv501(conv[501]),.conv502(conv[502]),.conv503(conv[503]),.conv504(conv[504]),.conv505(conv[505]),.conv506(conv[506]),.conv507(conv[507]),.conv508(conv[508]),.conv509(conv[509]),.conv510(conv[510]),.conv511(conv[511]),.conv512(conv[512]),.conv513(conv[513]),.conv514(conv[514]),.conv515(conv[515]),.conv516(conv[516]),.conv517(conv[517]),.conv518(conv[518]),.conv519(conv[519]),.conv520(conv[520]),.conv521(conv[521]),.conv522(conv[522]),.conv523(conv[523]),.conv524(conv[524]),.conv525(conv[525]),.conv526(conv[526]),.conv527(conv[527]),.conv528(conv[528]),.conv529(conv[529]),.conv530(conv[530]),.conv531(conv[531]),.conv532(conv[532]),.conv533(conv[533]),.conv534(conv[534]),.conv535(conv[535]),.conv536(conv[536]),.conv537(conv[537]),.conv538(conv[538]),.conv539(conv[539]),.conv540(conv[540]),.conv541(conv[541]),.conv542(conv[542]),.conv543(conv[543]),.conv544(conv[544]),.conv545(conv[545]),.conv546(conv[546]),.conv547(conv[547]),.conv548(conv[548]),.conv549(conv[549]),.conv550(conv[550]),.conv551(conv[551]),.conv552(conv[552]),.conv553(conv[553]),.conv554(conv[554]),.conv555(conv[555]),.conv556(conv[556]),.conv557(conv[557]),.conv558(conv[558]),.conv559(conv[559]),.conv560(conv[560]),.conv561(conv[561]),.conv562(conv[562]),.conv563(conv[563]),.conv564(conv[564]),.conv565(conv[565]),.conv566(conv[566]),.conv567(conv[567]),.conv568(conv[568]),.conv569(conv[569]),.conv570(conv[570]),.conv571(conv[571]),.conv572(conv[572]),.conv573(conv[573]),.conv574(conv[574]),.conv575(conv[575]),
.start(start));*/

/*FullyConnected FullyConnected1(.weight0(weight[0]),.weight1(weight[1]),.weight2(weight[2]),.weight3(weight[3]),.weight4(weight[4]),.weight5(weight[5]),.weight6(weight[6]),.weight7(weight[7]),.weight8(weight[8]),.weight9(weight[9]),.weight10(weight[10]),.weight11(weight[11]),.weight12(weight[12]),.weight13(weight[13]),.weight14(weight[14]),.weight15(weight[15]),.weight16(weight[16]),.weight17(weight[17]),.weight18(weight[18]),.weight19(weight[19]),.weight20(weight[20]),.weight21(weight[21]),.weight22(weight[22]),.weight23(weight[23]),.weight24(weight[24]),.weight25(weight[25]),.weight26(weight[26]),.weight27(weight[27]),.weight28(weight[28]),.weight29(weight[29]),.weight30(weight[30]),.weight31(weight[31]),.weight32(weight[32]),.weight33(weight[33]),.weight34(weight[34]),.weight35(weight[35]),.weight36(weight[36]),.weight37(weight[37]),.weight38(weight[38]),.weight39(weight[39]),.weight40(weight[40]),.weight41(weight[41]),.weight42(weight[42]),.weight43(weight[43]),.weight44(weight[44]),.weight45(weight[45]),.weight46(weight[46]),.weight47(weight[47]),.weight48(weight[48]),.weight49(weight[49]),.weight50(weight[50]),.weight51(weight[51]),.weight52(weight[52]),.weight53(weight[53]),.weight54(weight[54]),.weight55(weight[55]),.weight56(weight[56]),.weight57(weight[57]),.weight58(weight[58]),.weight59(weight[59]),.weight60(weight[60]),.weight61(weight[61]),.weight62(weight[62]),.weight63(weight[63]),.weight64(weight[64]),.weight65(weight[65]),.weight66(weight[66]),.weight67(weight[67]),.weight68(weight[68]),.weight69(weight[69]),.weight70(weight[70]),.weight71(weight[71]),.weight72(weight[72]),.weight73(weight[73]),.weight74(weight[74]),.weight75(weight[75]),.weight76(weight[76]),.weight77(weight[77]),.weight78(weight[78]),.weight79(weight[79]),.weight80(weight[80]),.weight81(weight[81]),.weight82(weight[82]),.weight83(weight[83]),.weight84(weight[84]),.weight85(weight[85]),.weight86(weight[86]),.weight87(weight[87]),.weight88(weight[88]),.weight89(weight[89]),.weight90(weight[90]),.weight91(weight[91]),.weight92(weight[92]),.weight93(weight[93]),.weight94(weight[94]),.weight95(weight[95]),.weight96(weight[96]),.weight97(weight[97]),.weight98(weight[98]),.weight99(weight[99]),.weight100(weight[100]),.weight101(weight[101]),.weight102(weight[102]),.weight103(weight[103]),.weight104(weight[104]),.weight105(weight[105]),.weight106(weight[106]),.weight107(weight[107]),.weight108(weight[108]),.weight109(weight[109]),.weight110(weight[110]),.weight111(weight[111]),.weight112(weight[112]),.weight113(weight[113]),.weight114(weight[114]),.weight115(weight[115]),.weight116(weight[116]),.weight117(weight[117]),.weight118(weight[118]),.weight119(weight[119]),.weight120(weight[120]),.weight121(weight[121]),.weight122(weight[122]),.weight123(weight[123]),.weight124(weight[124]),.weight125(weight[125]),.weight126(weight[126]),.weight127(weight[127]),.weight128(weight[128]),.weight129(weight[129]),.weight130(weight[130]),.weight131(weight[131]),.weight132(weight[132]),.weight133(weight[133]),.weight134(weight[134]),.weight135(weight[135]),.weight136(weight[136]),.weight137(weight[137]),.weight138(weight[138]),.weight139(weight[139]),.weight140(weight[140]),.weight141(weight[141]),.weight142(weight[142]),.weight143(weight[143]), .in0(in[0]),.in1(in[1]),.in2(in[2]),.in3(in[3]),.in4(in[4]),.in5(in[5]),.in6(in[6]),.in7(in[7]),.in8(in[8]),.in9(in[9]),.in10(in[10]),.in11(in[11]),.in12(in[12]),.in13(in[13]),.in14(in[14]),.in15(in[15]),.in16(in[16]),.in17(in[17]),.in18(in[18]),.in19(in[19]),.in20(in[20]),.in21(in[21]),.in22(in[22]),.in23(in[23]),.in24(in[24]),.in25(in[25]),.in26(in[26]),.in27(in[27]),.in28(in[28]),.in29(in[29]),.in30(in[30]),.in31(in[31]),.in32(in[32]),.in33(in[33]),.in34(in[34]),.in35(in[35]),.in36(in[36]),.in37(in[37]),.in38(in[38]),.in39(in[39]),.in40(in[40]),.in41(in[41]),.in42(in[42]),.in43(in[43]),.in44(in[44]),.in45(in[45]),.in46(in[46]),.in47(in[47]),.in48(in[48]),.in49(in[49]),.in50(in[50]),.in51(in[51]),.in52(in[52]),.in53(in[53]),.in54(in[54]),.in55(in[55]),.in56(in[56]),.in57(in[57]),.in58(in[58]),.in59(in[59]),.in60(in[60]),.in61(in[61]),.in62(in[62]),.in63(in[63]),.in64(in[64]),.in65(in[65]),.in66(in[66]),.in67(in[67]),.in68(in[68]),.in69(in[69]),.in70(in[70]),.in71(in[71]),.in72(in[72]),.in73(in[73]),.in74(in[74]),.in75(in[75]),.in76(in[76]),.in77(in[77]),.in78(in[78]),.in79(in[79]),.in80(in[80]),.in81(in[81]),.in82(in[82]),.in83(in[83]),.in84(in[84]),.in85(in[85]),.in86(in[86]),.in87(in[87]),.in88(in[88]),.in89(in[89]),.in90(in[90]),.in91(in[91]),.in92(in[92]),.in93(in[93]),.in94(in[94]),.in95(in[95]),.in96(in[96]),.in97(in[97]),.in98(in[98]),.in99(in[99]),.in100(in[100]),.in101(in[101]),.in102(in[102]),.in103(in[103]),.in104(in[104]),.in105(in[105]),.in106(in[106]),.in107(in[107]),.in108(in[108]),.in109(in[109]),.in110(in[110]),.in111(in[111]),.in112(in[112]),.in113(in[113]),.in114(in[114]),.in115(in[115]),.in116(in[116]),.in117(in[117]),.in118(in[118]),.in119(in[119]),.in120(in[120]),.in121(in[121]),.in122(in[122]),.in123(in[123]),.in124(in[124]),.in125(in[125]),.in126(in[126]),.in127(in[127]),.in128(in[128]),.in129(in[129]),.in130(in[130]),.in131(in[131]),.in132(in[132]),.in133(in[133]),.in134(in[134]),.in135(in[135]),.in136(in[136]),.in137(in[137]),.in138(in[138]),.in139(in[139]),.in140(in[140]),.in141(in[141]),.in142(in[142]),.in143(in[143]),.out(out),.clk(clk),.ready(ready),
.start(start));*/

always 
begin
#5 clk = !clk;
end


endmodule
